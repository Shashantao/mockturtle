module multiplier(q, a, b);
  wire _0000_;
  wire _0001_;
  wire _0002_;
  wire _0003_;
  wire _0004_;
  wire _0005_;
  wire _0006_;
  wire _0007_;
  wire _0008_;
  wire _0009_;
  wire _0010_;
  wire _0011_;
  wire _0012_;
  wire _0013_;
  wire _0014_;
  wire _0015_;
  wire _0016_;
  wire _0017_;
  wire _0018_;
  wire _0019_;
  wire _0020_;
  wire _0021_;
  wire _0022_;
  wire _0023_;
  wire _0024_;
  wire _0025_;
  wire _0026_;
  wire _0027_;
  wire _0028_;
  wire _0029_;
  wire _0030_;
  wire _0031_;
  wire _0032_;
  wire _0033_;
  wire _0034_;
  wire _0035_;
  wire _0036_;
  wire _0037_;
  wire _0038_;
  wire _0039_;
  wire _0040_;
  wire _0041_;
  wire _0042_;
  wire _0043_;
  wire _0044_;
  wire _0045_;
  wire _0046_;
  wire _0047_;
  wire _0048_;
  wire _0049_;
  wire _0050_;
  wire _0051_;
  wire _0052_;
  wire _0053_;
  wire _0054_;
  wire _0055_;
  wire _0056_;
  wire _0057_;
  wire _0058_;
  wire _0059_;
  wire _0060_;
  wire _0061_;
  wire _0062_;
  wire _0063_;
  wire _0064_;
  wire _0065_;
  wire _0066_;
  wire _0067_;
  wire _0068_;
  wire _0069_;
  wire _0070_;
  wire _0071_;
  wire _0072_;
  wire _0073_;
  wire _0074_;
  wire _0075_;
  wire _0076_;
  wire _0077_;
  wire _0078_;
  wire _0079_;
  wire _0080_;
  wire _0081_;
  wire _0082_;
  wire _0083_;
  wire _0084_;
  wire _0085_;
  wire _0086_;
  wire _0087_;
  wire _0088_;
  wire _0089_;
  wire _0090_;
  wire _0091_;
  wire _0092_;
  wire _0093_;
  wire _0094_;
  wire _0095_;
  wire _0096_;
  wire _0097_;
  wire _0098_;
  wire _0099_;
  wire _0100_;
  wire _0101_;
  wire _0102_;
  wire _0103_;
  wire _0104_;
  wire _0105_;
  wire _0106_;
  wire _0107_;
  wire _0108_;
  wire _0109_;
  wire _0110_;
  wire _0111_;
  wire _0112_;
  wire _0113_;
  wire _0114_;
  wire _0115_;
  wire _0116_;
  wire _0117_;
  wire _0118_;
  wire _0119_;
  wire _0120_;
  wire _0121_;
  wire _0122_;
  wire _0123_;
  wire _0124_;
  wire _0125_;
  wire _0126_;
  wire _0127_;
  wire _0128_;
  wire _0129_;
  wire _0130_;
  wire _0131_;
  wire _0132_;
  wire _0133_;
  wire _0134_;
  wire _0135_;
  wire _0136_;
  wire _0137_;
  wire _0138_;
  wire _0139_;
  wire _0140_;
  wire _0141_;
  wire _0142_;
  wire _0143_;
  wire _0144_;
  wire _0145_;
  wire _0146_;
  wire _0147_;
  wire _0148_;
  wire _0149_;
  wire _0150_;
  wire _0151_;
  wire _0152_;
  wire _0153_;
  wire _0154_;
  wire _0155_;
  wire _0156_;
  wire _0157_;
  wire _0158_;
  wire _0159_;
  wire _0160_;
  wire _0161_;
  wire _0162_;
  wire _0163_;
  wire _0164_;
  wire _0165_;
  wire _0166_;
  wire _0167_;
  wire _0168_;
  wire _0169_;
  wire _0170_;
  wire _0171_;
  wire _0172_;
  wire _0173_;
  wire _0174_;
  wire _0175_;
  wire _0176_;
  wire _0177_;
  wire _0178_;
  wire _0179_;
  wire _0180_;
  wire _0181_;
  wire _0182_;
  wire _0183_;
  wire _0184_;
  wire _0185_;
  wire _0186_;
  wire _0187_;
  wire _0188_;
  wire _0189_;
  wire _0190_;
  wire _0191_;
  wire _0192_;
  wire _0193_;
  wire _0194_;
  wire _0195_;
  wire _0196_;
  wire _0197_;
  wire _0198_;
  wire _0199_;
  wire _0200_;
  wire _0201_;
  wire _0202_;
  wire _0203_;
  wire _0204_;
  wire _0205_;
  wire _0206_;
  wire _0207_;
  wire _0208_;
  wire _0209_;
  wire _0210_;
  wire _0211_;
  wire _0212_;
  wire _0213_;
  wire _0214_;
  wire _0215_;
  wire _0216_;
  wire _0217_;
  wire _0218_;
  wire _0219_;
  wire _0220_;
  wire _0221_;
  wire _0222_;
  wire _0223_;
  wire _0224_;
  wire _0225_;
  wire _0226_;
  wire _0227_;
  wire _0228_;
  wire _0229_;
  wire _0230_;
  wire _0231_;
  wire _0232_;
  wire _0233_;
  wire _0234_;
  wire _0235_;
  wire _0236_;
  wire _0237_;
  wire _0238_;
  wire _0239_;
  wire _0240_;
  wire _0241_;
  wire _0242_;
  wire _0243_;
  wire _0244_;
  wire _0245_;
  wire _0246_;
  wire _0247_;
  wire _0248_;
  wire _0249_;
  wire _0250_;
  wire _0251_;
  wire _0252_;
  wire _0253_;
  wire _0254_;
  wire _0255_;
  wire _0256_;
  wire _0257_;
  wire _0258_;
  wire _0259_;
  wire _0260_;
  wire _0261_;
  wire _0262_;
  wire _0263_;
  wire _0264_;
  wire _0265_;
  wire _0266_;
  wire _0267_;
  wire _0268_;
  wire _0269_;
  wire _0270_;
  wire _0271_;
  wire _0272_;
  wire _0273_;
  wire _0274_;
  wire _0275_;
  wire _0276_;
  wire _0277_;
  wire _0278_;
  wire _0279_;
  wire _0280_;
  wire _0281_;
  wire _0282_;
  wire _0283_;
  wire _0284_;
  wire _0285_;
  wire _0286_;
  wire _0287_;
  wire _0288_;
  wire _0289_;
  wire _0290_;
  wire _0291_;
  wire _0292_;
  wire _0293_;
  wire _0294_;
  wire _0295_;
  wire _0296_;
  wire _0297_;
  wire _0298_;
  wire _0299_;
  wire _0300_;
  wire _0301_;
  wire _0302_;
  wire _0303_;
  wire _0304_;
  wire _0305_;
  wire _0306_;
  wire _0307_;
  wire _0308_;
  wire _0309_;
  wire _0310_;
  wire _0311_;
  wire _0312_;
  wire _0313_;
  wire _0314_;
  wire _0315_;
  wire _0316_;
  wire _0317_;
  wire _0318_;
  wire _0319_;
  wire _0320_;
  wire _0321_;
  wire _0322_;
  wire _0323_;
  wire _0324_;
  wire _0325_;
  wire _0326_;
  wire _0327_;
  wire _0328_;
  wire _0329_;
  wire _0330_;
  wire _0331_;
  wire _0332_;
  wire _0333_;
  wire _0334_;
  wire _0335_;
  wire _0336_;
  wire _0337_;
  wire _0338_;
  wire _0339_;
  wire _0340_;
  wire _0341_;
  wire _0342_;
  wire _0343_;
  wire _0344_;
  wire _0345_;
  wire _0346_;
  wire _0347_;
  wire _0348_;
  wire _0349_;
  wire _0350_;
  wire _0351_;
  wire _0352_;
  wire _0353_;
  wire _0354_;
  wire _0355_;
  wire _0356_;
  wire _0357_;
  wire _0358_;
  wire _0359_;
  wire _0360_;
  wire _0361_;
  wire _0362_;
  wire _0363_;
  wire _0364_;
  wire _0365_;
  wire _0366_;
  wire _0367_;
  wire _0368_;
  wire _0369_;
  wire _0370_;
  wire _0371_;
  wire _0372_;
  wire _0373_;
  wire _0374_;
  wire _0375_;
  wire _0376_;
  wire _0377_;
  wire _0378_;
  wire _0379_;
  wire _0380_;
  wire _0381_;
  wire _0382_;
  wire _0383_;
  wire _0384_;
  wire _0385_;
  wire _0386_;
  wire _0387_;
  wire _0388_;
  wire _0389_;
  wire _0390_;
  wire _0391_;
  wire _0392_;
  wire _0393_;
  wire _0394_;
  wire _0395_;
  wire _0396_;
  wire _0397_;
  wire _0398_;
  wire _0399_;
  wire _0400_;
  wire _0401_;
  wire _0402_;
  wire _0403_;
  wire _0404_;
  wire _0405_;
  wire _0406_;
  wire _0407_;
  wire _0408_;
  wire _0409_;
  wire _0410_;
  wire _0411_;
  wire _0412_;
  wire _0413_;
  wire _0414_;
  wire _0415_;
  wire _0416_;
  wire _0417_;
  wire _0418_;
  wire _0419_;
  wire _0420_;
  wire _0421_;
  wire _0422_;
  wire _0423_;
  wire _0424_;
  wire _0425_;
  wire _0426_;
  wire _0427_;
  wire _0428_;
  wire _0429_;
  wire _0430_;
  wire _0431_;
  wire _0432_;
  wire _0433_;
  wire _0434_;
  wire _0435_;
  wire _0436_;
  wire _0437_;
  wire _0438_;
  wire _0439_;
  wire _0440_;
  wire _0441_;
  wire _0442_;
  wire _0443_;
  wire _0444_;
  wire _0445_;
  wire _0446_;
  wire _0447_;
  wire _0448_;
  wire _0449_;
  wire _0450_;
  wire _0451_;
  wire _0452_;
  wire _0453_;
  wire _0454_;
  wire _0455_;
  wire _0456_;
  wire _0457_;
  wire _0458_;
  wire _0459_;
  wire _0460_;
  wire _0461_;
  wire _0462_;
  wire _0463_;
  wire _0464_;
  wire _0465_;
  wire _0466_;
  wire _0467_;
  wire _0468_;
  wire _0469_;
  wire _0470_;
  wire _0471_;
  wire _0472_;
  wire _0473_;
  wire _0474_;
  wire _0475_;
  wire _0476_;
  wire _0477_;
  wire _0478_;
  wire _0479_;
  wire _0480_;
  wire _0481_;
  wire _0482_;
  wire _0483_;
  wire _0484_;
  wire _0485_;
  wire _0486_;
  wire _0487_;
  wire _0488_;
  wire _0489_;
  wire _0490_;
  wire _0491_;
  wire _0492_;
  wire _0493_;
  wire _0494_;
  wire _0495_;
  wire _0496_;
  wire _0497_;
  wire _0498_;
  wire _0499_;
  wire _0500_;
  wire _0501_;
  wire _0502_;
  wire _0503_;
  wire _0504_;
  wire _0505_;
  wire _0506_;
  wire _0507_;
  wire _0508_;
  wire _0509_;
  wire _0510_;
  wire _0511_;
  wire _0512_;
  wire _0513_;
  wire _0514_;
  wire _0515_;
  wire _0516_;
  wire _0517_;
  wire _0518_;
  wire _0519_;
  wire _0520_;
  wire _0521_;
  wire _0522_;
  wire _0523_;
  wire _0524_;
  wire _0525_;
  wire _0526_;
  wire _0527_;
  wire _0528_;
  wire _0529_;
  wire _0530_;
  wire _0531_;
  wire _0532_;
  wire _0533_;
  wire _0534_;
  wire _0535_;
  wire _0536_;
  wire _0537_;
  wire _0538_;
  wire _0539_;
  wire _0540_;
  wire _0541_;
  wire _0542_;
  wire _0543_;
  wire _0544_;
  wire _0545_;
  wire _0546_;
  wire _0547_;
  wire _0548_;
  wire _0549_;
  wire _0550_;
  wire _0551_;
  wire _0552_;
  wire _0553_;
  wire _0554_;
  wire _0555_;
  wire _0556_;
  wire _0557_;
  wire _0558_;
  wire _0559_;
  wire _0560_;
  wire _0561_;
  wire _0562_;
  wire _0563_;
  wire _0564_;
  wire _0565_;
  wire _0566_;
  wire _0567_;
  wire _0568_;
  wire _0569_;
  wire _0570_;
  wire _0571_;
  wire _0572_;
  wire _0573_;
  wire _0574_;
  wire _0575_;
  wire _0576_;
  wire _0577_;
  wire _0578_;
  wire _0579_;
  wire _0580_;
  wire _0581_;
  wire _0582_;
  wire _0583_;
  wire _0584_;
  wire _0585_;
  wire _0586_;
  wire _0587_;
  wire _0588_;
  wire _0589_;
  wire _0590_;
  wire _0591_;
  wire _0592_;
  wire _0593_;
  wire _0594_;
  wire _0595_;
  wire _0596_;
  wire _0597_;
  wire _0598_;
  wire _0599_;
  wire _0600_;
  wire _0601_;
  wire _0602_;
  wire _0603_;
  wire _0604_;
  wire _0605_;
  wire _0606_;
  wire _0607_;
  wire _0608_;
  wire _0609_;
  wire _0610_;
  wire _0611_;
  wire _0612_;
  wire _0613_;
  wire _0614_;
  wire _0615_;
  wire _0616_;
  wire _0617_;
  wire _0618_;
  wire _0619_;
  wire _0620_;
  wire _0621_;
  wire _0622_;
  wire _0623_;
  wire _0624_;
  wire _0625_;
  wire _0626_;
  wire _0627_;
  wire _0628_;
  wire _0629_;
  wire _0630_;
  wire _0631_;
  wire _0632_;
  wire _0633_;
  wire _0634_;
  wire _0635_;
  wire _0636_;
  wire _0637_;
  wire _0638_;
  wire _0639_;
  wire _0640_;
  wire _0641_;
  wire _0642_;
  wire _0643_;
  wire _0644_;
  wire _0645_;
  wire _0646_;
  wire _0647_;
  wire _0648_;
  wire _0649_;
  wire _0650_;
  wire _0651_;
  wire _0652_;
  wire _0653_;
  wire _0654_;
  wire _0655_;
  wire _0656_;
  wire _0657_;
  wire _0658_;
  wire _0659_;
  wire _0660_;
  wire _0661_;
  wire _0662_;
  wire _0663_;
  wire _0664_;
  wire _0665_;
  wire _0666_;
  wire _0667_;
  wire _0668_;
  wire _0669_;
  wire _0670_;
  wire _0671_;
  wire _0672_;
  wire _0673_;
  wire _0674_;
  wire _0675_;
  wire _0676_;
  wire _0677_;
  wire _0678_;
  wire _0679_;
  wire _0680_;
  wire _0681_;
  wire _0682_;
  wire _0683_;
  wire _0684_;
  wire _0685_;
  wire _0686_;
  wire _0687_;
  wire _0688_;
  wire _0689_;
  wire _0690_;
  wire _0691_;
  wire _0692_;
  wire _0693_;
  wire _0694_;
  wire _0695_;
  wire _0696_;
  wire _0697_;
  wire _0698_;
  wire _0699_;
  wire _0700_;
  wire _0701_;
  wire _0702_;
  wire _0703_;
  wire _0704_;
  wire _0705_;
  wire _0706_;
  wire _0707_;
  wire _0708_;
  wire _0709_;
  wire _0710_;
  wire _0711_;
  wire _0712_;
  wire _0713_;
  wire _0714_;
  wire _0715_;
  wire _0716_;
  wire _0717_;
  wire _0718_;
  wire _0719_;
  wire _0720_;
  wire _0721_;
  wire _0722_;
  wire _0723_;
  wire _0724_;
  wire _0725_;
  wire _0726_;
  wire _0727_;
  wire _0728_;
  wire _0729_;
  wire _0730_;
  wire _0731_;
  wire _0732_;
  wire _0733_;
  wire _0734_;
  wire _0735_;
  wire _0736_;
  wire _0737_;
  wire _0738_;
  wire _0739_;
  wire _0740_;
  wire _0741_;
  wire _0742_;
  wire _0743_;
  wire _0744_;
  wire _0745_;
  wire _0746_;
  wire _0747_;
  wire _0748_;
  wire _0749_;
  wire _0750_;
  wire _0751_;
  wire _0752_;
  wire _0753_;
  wire _0754_;
  wire _0755_;
  wire _0756_;
  wire _0757_;
  wire _0758_;
  wire _0759_;
  wire _0760_;
  wire _0761_;
  wire _0762_;
  wire _0763_;
  wire _0764_;
  wire _0765_;
  wire _0766_;
  wire _0767_;
  wire _0768_;
  wire _0769_;
  wire _0770_;
  wire _0771_;
  wire _0772_;
  wire _0773_;
  wire _0774_;
  wire _0775_;
  wire _0776_;
  wire _0777_;
  wire _0778_;
  wire _0779_;
  wire _0780_;
  wire _0781_;
  wire _0782_;
  wire _0783_;
  wire _0784_;
  wire _0785_;
  wire _0786_;
  wire _0787_;
  wire _0788_;
  wire _0789_;
  wire _0790_;
  wire _0791_;
  wire _0792_;
  wire _0793_;
  wire _0794_;
  wire _0795_;
  wire _0796_;
  wire _0797_;
  wire _0798_;
  wire _0799_;
  wire _0800_;
  wire _0801_;
  wire _0802_;
  wire _0803_;
  wire _0804_;
  wire _0805_;
  wire _0806_;
  wire _0807_;
  wire _0808_;
  wire _0809_;
  wire _0810_;
  wire _0811_;
  wire _0812_;
  wire _0813_;
  wire _0814_;
  wire _0815_;
  wire _0816_;
  wire _0817_;
  wire _0818_;
  wire _0819_;
  wire _0820_;
  wire _0821_;
  wire _0822_;
  wire _0823_;
  wire _0824_;
  wire _0825_;
  wire _0826_;
  wire _0827_;
  wire _0828_;
  wire _0829_;
  wire _0830_;
  wire _0831_;
  wire _0832_;
  wire _0833_;
  wire _0834_;
  wire _0835_;
  wire _0836_;
  wire _0837_;
  wire _0838_;
  wire _0839_;
  wire _0840_;
  wire _0841_;
  wire _0842_;
  wire _0843_;
  wire _0844_;
  wire _0845_;
  wire _0846_;
  wire _0847_;
  wire _0848_;
  wire _0849_;
  wire _0850_;
  wire _0851_;
  wire _0852_;
  wire _0853_;
  wire _0854_;
  wire _0855_;
  wire _0856_;
  wire _0857_;
  wire _0858_;
  wire _0859_;
  wire _0860_;
  wire _0861_;
  wire _0862_;
  wire _0863_;
  wire _0864_;
  wire _0865_;
  wire _0866_;
  wire _0867_;
  wire _0868_;
  wire _0869_;
  wire _0870_;
  wire _0871_;
  wire _0872_;
  wire _0873_;
  wire _0874_;
  wire _0875_;
  wire _0876_;
  wire _0877_;
  wire _0878_;
  wire _0879_;
  wire _0880_;
  wire _0881_;
  wire _0882_;
  wire _0883_;
  wire _0884_;
  wire _0885_;
  wire _0886_;
  wire _0887_;
  wire _0888_;
  wire _0889_;
  wire _0890_;
  wire _0891_;
  wire _0892_;
  wire _0893_;
  wire _0894_;
  wire _0895_;
  wire _0896_;
  wire _0897_;
  wire _0898_;
  wire _0899_;
  wire _0900_;
  wire _0901_;
  wire _0902_;
  wire _0903_;
  wire _0904_;
  wire _0905_;
  wire _0906_;
  wire _0907_;
  wire _0908_;
  wire _0909_;
  wire _0910_;
  wire _0911_;
  wire _0912_;
  wire _0913_;
  wire _0914_;
  wire _0915_;
  wire _0916_;
  wire _0917_;
  wire _0918_;
  wire _0919_;
  wire _0920_;
  wire _0921_;
  wire _0922_;
  wire _0923_;
  wire _0924_;
  wire _0925_;
  wire _0926_;
  wire _0927_;
  wire _0928_;
  wire _0929_;
  wire _0930_;
  wire _0931_;
  wire _0932_;
  wire _0933_;
  wire _0934_;
  wire _0935_;
  wire _0936_;
  wire _0937_;
  wire _0938_;
  wire _0939_;
  wire _0940_;
  wire _0941_;
  wire _0942_;
  wire _0943_;
  wire _0944_;
  wire _0945_;
  wire _0946_;
  wire _0947_;
  wire _0948_;
  wire _0949_;
  wire _0950_;
  wire _0951_;
  wire _0952_;
  wire _0953_;
  wire _0954_;
  wire _0955_;
  wire _0956_;
  wire _0957_;
  wire _0958_;
  wire _0959_;
  wire _0960_;
  wire _0961_;
  wire _0962_;
  wire _0963_;
  wire _0964_;
  wire _0965_;
  wire _0966_;
  wire _0967_;
  wire _0968_;
  wire _0969_;
  wire _0970_;
  wire _0971_;
  wire _0972_;
  wire _0973_;
  wire _0974_;
  wire _0975_;
  wire _0976_;
  wire _0977_;
  wire _0978_;
  wire _0979_;
  wire _0980_;
  wire _0981_;
  wire _0982_;
  wire _0983_;
  wire _0984_;
  wire _0985_;
  wire _0986_;
  wire _0987_;
  wire _0988_;
  wire _0989_;
  wire _0990_;
  wire _0991_;
  wire _0992_;
  wire _0993_;
  wire _0994_;
  wire _0995_;
  wire _0996_;
  wire _0997_;
  wire _0998_;
  wire _0999_;
  wire _1000_;
  wire _1001_;
  wire _1002_;
  wire _1003_;
  wire _1004_;
  wire _1005_;
  wire _1006_;
  wire _1007_;
  wire _1008_;
  wire _1009_;
  wire _1010_;
  wire _1011_;
  wire _1012_;
  wire _1013_;
  wire _1014_;
  wire _1015_;
  wire _1016_;
  wire _1017_;
  wire _1018_;
  wire _1019_;
  wire _1020_;
  wire _1021_;
  wire _1022_;
  wire _1023_;
  wire _1024_;
  wire _1025_;
  wire _1026_;
  wire _1027_;
  wire _1028_;
  wire _1029_;
  wire _1030_;
  wire _1031_;
  wire _1032_;
  wire _1033_;
  wire _1034_;
  wire _1035_;
  wire _1036_;
  wire _1037_;
  wire _1038_;
  wire _1039_;
  wire _1040_;
  wire _1041_;
  wire _1042_;
  wire _1043_;
  wire _1044_;
  wire _1045_;
  wire _1046_;
  wire _1047_;
  wire _1048_;
  wire _1049_;
  wire _1050_;
  wire _1051_;
  wire _1052_;
  wire _1053_;
  wire _1054_;
  wire _1055_;
  wire _1056_;
  wire _1057_;
  wire _1058_;
  wire _1059_;
  wire _1060_;
  wire _1061_;
  wire _1062_;
  wire _1063_;
  wire _1064_;
  wire _1065_;
  wire _1066_;
  wire _1067_;
  wire _1068_;
  wire _1069_;
  wire _1070_;
  wire _1071_;
  wire _1072_;
  wire _1073_;
  wire _1074_;
  wire _1075_;
  wire _1076_;
  wire _1077_;
  wire _1078_;
  wire _1079_;
  wire _1080_;
  wire _1081_;
  wire _1082_;
  wire _1083_;
  wire _1084_;
  wire _1085_;
  wire _1086_;
  wire _1087_;
  wire _1088_;
  wire _1089_;
  wire _1090_;
  wire _1091_;
  wire _1092_;
  wire _1093_;
  wire _1094_;
  wire _1095_;
  wire _1096_;
  wire _1097_;
  wire _1098_;
  wire _1099_;
  wire _1100_;
  wire _1101_;
  wire _1102_;
  wire _1103_;
  wire _1104_;
  wire _1105_;
  wire _1106_;
  wire _1107_;
  wire _1108_;
  wire _1109_;
  wire _1110_;
  wire _1111_;
  wire _1112_;
  wire _1113_;
  wire _1114_;
  wire _1115_;
  wire _1116_;
  wire _1117_;
  wire _1118_;
  wire _1119_;
  wire _1120_;
  wire _1121_;
  wire _1122_;
  wire _1123_;
  wire _1124_;
  wire _1125_;
  wire _1126_;
  wire _1127_;
  wire _1128_;
  wire _1129_;
  wire _1130_;
  wire _1131_;
  wire _1132_;
  wire _1133_;
  wire _1134_;
  wire _1135_;
  wire _1136_;
  wire _1137_;
  wire _1138_;
  wire _1139_;
  wire _1140_;
  wire _1141_;
  wire _1142_;
  wire _1143_;
  wire _1144_;
  wire _1145_;
  wire _1146_;
  wire _1147_;
  wire _1148_;
  wire _1149_;
  wire _1150_;
  wire _1151_;
  wire _1152_;
  wire _1153_;
  wire _1154_;
  wire _1155_;
  wire _1156_;
  wire _1157_;
  wire _1158_;
  wire _1159_;
  wire _1160_;
  wire _1161_;
  wire _1162_;
  wire _1163_;
  wire _1164_;
  wire _1165_;
  wire _1166_;
  wire _1167_;
  wire _1168_;
  wire _1169_;
  wire _1170_;
  wire _1171_;
  wire _1172_;
  wire _1173_;
  wire _1174_;
  wire _1175_;
  wire _1176_;
  wire _1177_;
  wire _1178_;
  wire _1179_;
  wire _1180_;
  wire _1181_;
  wire _1182_;
  wire _1183_;
  wire _1184_;
  wire _1185_;
  wire _1186_;
  wire _1187_;
  wire _1188_;
  wire _1189_;
  wire _1190_;
  wire _1191_;
  wire _1192_;
  wire _1193_;
  wire _1194_;
  wire _1195_;
  wire _1196_;
  wire _1197_;
  wire _1198_;
  wire _1199_;
  wire _1200_;
  wire _1201_;
  wire _1202_;
  wire _1203_;
  wire _1204_;
  wire _1205_;
  wire _1206_;
  wire _1207_;
  wire _1208_;
  wire _1209_;
  wire _1210_;
  wire _1211_;
  wire _1212_;
  wire _1213_;
  wire _1214_;
  wire _1215_;
  wire _1216_;
  wire _1217_;
  wire _1218_;
  wire _1219_;
  wire _1220_;
  wire _1221_;
  wire _1222_;
  wire _1223_;
  wire _1224_;
  wire _1225_;
  wire _1226_;
  wire _1227_;
  wire _1228_;
  wire _1229_;
  wire _1230_;
  wire _1231_;
  wire _1232_;
  wire _1233_;
  wire _1234_;
  wire _1235_;
  wire _1236_;
  wire _1237_;
  wire _1238_;
  wire _1239_;
  wire _1240_;
  wire _1241_;
  wire _1242_;
  wire _1243_;
  wire _1244_;
  wire _1245_;
  wire _1246_;
  wire _1247_;
  wire _1248_;
  wire _1249_;
  wire _1250_;
  wire _1251_;
  wire _1252_;
  wire _1253_;
  wire _1254_;
  wire _1255_;
  wire _1256_;
  wire _1257_;
  wire _1258_;
  wire _1259_;
  wire _1260_;
  wire _1261_;
  wire _1262_;
  wire _1263_;
  wire _1264_;
  wire _1265_;
  wire _1266_;
  wire _1267_;
  wire _1268_;
  wire _1269_;
  wire _1270_;
  wire _1271_;
  wire _1272_;
  wire _1273_;
  wire _1274_;
  wire _1275_;
  wire _1276_;
  wire _1277_;
  wire _1278_;
  wire _1279_;
  wire _1280_;
  wire _1281_;
  wire _1282_;
  wire _1283_;
  wire _1284_;
  wire _1285_;
  wire _1286_;
  wire _1287_;
  wire _1288_;
  wire _1289_;
  wire _1290_;
  wire _1291_;
  wire _1292_;
  wire _1293_;
  wire _1294_;
  wire _1295_;
  wire _1296_;
  wire _1297_;
  wire _1298_;
  wire _1299_;
  wire _1300_;
  wire _1301_;
  wire _1302_;
  wire _1303_;
  wire _1304_;
  wire _1305_;
  wire _1306_;
  wire _1307_;
  wire _1308_;
  wire _1309_;
  wire _1310_;
  wire _1311_;
  wire _1312_;
  wire _1313_;
  wire _1314_;
  wire _1315_;
  wire _1316_;
  wire _1317_;
  wire _1318_;
  wire _1319_;
  wire _1320_;
  wire _1321_;
  wire _1322_;
  wire _1323_;
  wire _1324_;
  wire _1325_;
  wire _1326_;
  wire _1327_;
  wire _1328_;
  wire _1329_;
  wire _1330_;
  wire _1331_;
  wire _1332_;
  wire _1333_;
  wire _1334_;
  wire _1335_;
  wire _1336_;
  wire _1337_;
  wire _1338_;
  wire _1339_;
  wire _1340_;
  wire _1341_;
  wire _1342_;
  wire _1343_;
  wire _1344_;
  wire _1345_;
  wire _1346_;
  wire _1347_;
  wire _1348_;
  wire _1349_;
  wire _1350_;
  wire _1351_;
  wire _1352_;
  wire _1353_;
  wire _1354_;
  wire _1355_;
  wire _1356_;
  wire _1357_;
  wire _1358_;
  wire _1359_;
  wire _1360_;
  wire _1361_;
  wire _1362_;
  wire _1363_;
  wire _1364_;
  wire _1365_;
  wire _1366_;
  wire _1367_;
  wire _1368_;
  wire _1369_;
  wire _1370_;
  wire _1371_;
  wire _1372_;
  wire _1373_;
  wire _1374_;
  wire _1375_;
  wire _1376_;
  wire _1377_;
  wire _1378_;
  wire _1379_;
  wire _1380_;
  wire _1381_;
  wire _1382_;
  wire _1383_;
  wire _1384_;
  wire _1385_;
  wire _1386_;
  wire _1387_;
  wire _1388_;
  wire _1389_;
  wire _1390_;
  wire _1391_;
  wire _1392_;
  wire _1393_;
  wire _1394_;
  wire _1395_;
  wire _1396_;
  wire _1397_;
  wire _1398_;
  wire _1399_;
  wire _1400_;
  wire _1401_;
  wire _1402_;
  wire _1403_;
  wire _1404_;
  wire _1405_;
  wire _1406_;
  wire _1407_;
  wire _1408_;
  wire _1409_;
  wire _1410_;
  wire _1411_;
  wire _1412_;
  wire _1413_;
  wire _1414_;
  wire _1415_;
  wire _1416_;
  wire _1417_;
  wire _1418_;
  wire _1419_;
  wire _1420_;
  wire _1421_;
  wire _1422_;
  wire _1423_;
  wire _1424_;
  wire _1425_;
  wire _1426_;
  wire _1427_;
  wire _1428_;
  wire _1429_;
  wire _1430_;
  wire _1431_;
  wire _1432_;
  wire _1433_;
  wire _1434_;
  wire _1435_;
  wire _1436_;
  wire _1437_;
  wire _1438_;
  wire _1439_;
  wire _1440_;
  wire _1441_;
  wire _1442_;
  wire _1443_;
  wire _1444_;
  wire _1445_;
  wire _1446_;
  wire _1447_;
  wire _1448_;
  wire _1449_;
  wire _1450_;
  wire _1451_;
  wire _1452_;
  wire _1453_;
  wire _1454_;
  wire _1455_;
  wire _1456_;
  wire _1457_;
  wire _1458_;
  wire _1459_;
  wire _1460_;
  wire _1461_;
  wire _1462_;
  wire _1463_;
  wire _1464_;
  wire _1465_;
  wire _1466_;
  wire _1467_;
  wire _1468_;
  wire _1469_;
  wire _1470_;
  wire _1471_;
  wire _1472_;
  wire _1473_;
  wire _1474_;
  wire _1475_;
  wire _1476_;
  wire _1477_;
  wire _1478_;
  wire _1479_;
  wire _1480_;
  wire _1481_;
  wire _1482_;
  wire _1483_;
  wire _1484_;
  wire _1485_;
  wire _1486_;
  wire _1487_;
  wire _1488_;
  wire _1489_;
  wire _1490_;
  wire _1491_;
  wire _1492_;
  wire _1493_;
  wire _1494_;
  wire _1495_;
  wire _1496_;
  wire _1497_;
  wire _1498_;
  wire _1499_;
  wire _1500_;
  wire _1501_;
  wire _1502_;
  wire _1503_;
  wire _1504_;
  wire _1505_;
  wire _1506_;
  wire _1507_;
  wire _1508_;
  wire _1509_;
  wire _1510_;
  wire _1511_;
  wire _1512_;
  wire _1513_;
  wire _1514_;
  wire _1515_;
  wire _1516_;
  wire _1517_;
  wire _1518_;
  wire _1519_;
  wire _1520_;
  wire _1521_;
  wire _1522_;
  wire _1523_;
  wire _1524_;
  wire _1525_;
  wire _1526_;
  wire _1527_;
  wire _1528_;
  wire _1529_;
  wire _1530_;
  wire _1531_;
  wire _1532_;
  wire _1533_;
  wire _1534_;
  wire _1535_;
  wire _1536_;
  wire _1537_;
  wire _1538_;
  wire _1539_;
  wire _1540_;
  wire _1541_;
  wire _1542_;
  wire _1543_;
  wire _1544_;
  wire _1545_;
  wire _1546_;
  wire _1547_;
  wire _1548_;
  wire _1549_;
  wire _1550_;
  wire _1551_;
  wire _1552_;
  wire _1553_;
  wire _1554_;
  wire _1555_;
  wire _1556_;
  wire _1557_;
  wire _1558_;
  wire _1559_;
  wire _1560_;
  wire _1561_;
  wire _1562_;
  wire _1563_;
  wire _1564_;
  wire _1565_;
  wire _1566_;
  wire _1567_;
  wire _1568_;
  wire _1569_;
  wire _1570_;
  wire _1571_;
  wire _1572_;
  wire _1573_;
  wire _1574_;
  wire _1575_;
  wire _1576_;
  wire _1577_;
  wire _1578_;
  wire _1579_;
  wire _1580_;
  wire _1581_;
  wire _1582_;
  wire _1583_;
  wire _1584_;
  wire _1585_;
  wire _1586_;
  wire _1587_;
  wire _1588_;
  wire _1589_;
  wire _1590_;
  wire _1591_;
  wire _1592_;
  wire _1593_;
  wire _1594_;
  wire _1595_;
  wire _1596_;
  wire _1597_;
  wire _1598_;
  wire _1599_;
  wire _1600_;
  wire _1601_;
  wire _1602_;
  wire _1603_;
  wire _1604_;
  wire _1605_;
  wire _1606_;
  wire _1607_;
  wire _1608_;
  wire _1609_;
  wire _1610_;
  wire _1611_;
  wire _1612_;
  wire _1613_;
  wire _1614_;
  wire _1615_;
  wire _1616_;
  wire _1617_;
  wire _1618_;
  wire _1619_;
  wire _1620_;
  wire _1621_;
  wire _1622_;
  wire _1623_;
  wire _1624_;
  wire _1625_;
  wire _1626_;
  wire _1627_;
  wire _1628_;
  wire _1629_;
  wire _1630_;
  wire _1631_;
  wire _1632_;
  wire _1633_;
  wire _1634_;
  wire _1635_;
  wire _1636_;
  wire _1637_;
  wire _1638_;
  wire _1639_;
  wire _1640_;
  wire _1641_;
  wire _1642_;
  wire _1643_;
  wire _1644_;
  wire _1645_;
  wire _1646_;
  wire _1647_;
  wire _1648_;
  wire _1649_;
  wire _1650_;
  wire _1651_;
  wire _1652_;
  wire _1653_;
  wire _1654_;
  wire _1655_;
  wire _1656_;
  wire _1657_;
  wire _1658_;
  wire _1659_;
  wire _1660_;
  wire _1661_;
  wire _1662_;
  wire _1663_;
  wire _1664_;
  wire _1665_;
  wire _1666_;
  wire _1667_;
  wire _1668_;
  wire _1669_;
  wire _1670_;
  wire _1671_;
  wire _1672_;
  wire _1673_;
  wire _1674_;
  wire _1675_;
  wire _1676_;
  wire _1677_;
  wire _1678_;
  wire _1679_;
  wire _1680_;
  wire _1681_;
  wire _1682_;
  wire _1683_;
  wire _1684_;
  wire _1685_;
  wire _1686_;
  wire _1687_;
  wire _1688_;
  wire _1689_;
  wire _1690_;
  wire _1691_;
  wire _1692_;
  wire _1693_;
  wire _1694_;
  wire _1695_;
  wire _1696_;
  wire _1697_;
  wire _1698_;
  wire _1699_;
  wire _1700_;
  wire _1701_;
  wire _1702_;
  wire _1703_;
  wire _1704_;
  wire _1705_;
  wire _1706_;
  wire _1707_;
  wire _1708_;
  wire _1709_;
  wire _1710_;
  wire _1711_;
  wire _1712_;
  wire _1713_;
  wire _1714_;
  wire _1715_;
  wire _1716_;
  wire _1717_;
  wire _1718_;
  wire _1719_;
  wire _1720_;
  wire _1721_;
  wire _1722_;
  wire _1723_;
  wire _1724_;
  wire _1725_;
  wire _1726_;
  wire _1727_;
  wire _1728_;
  wire _1729_;
  wire _1730_;
  wire _1731_;
  wire _1732_;
  wire _1733_;
  wire _1734_;
  wire _1735_;
  wire _1736_;
  wire _1737_;
  wire _1738_;
  wire _1739_;
  wire _1740_;
  wire _1741_;
  wire _1742_;
  wire _1743_;
  wire _1744_;
  wire _1745_;
  wire _1746_;
  wire _1747_;
  wire _1748_;
  wire _1749_;
  wire _1750_;
  wire _1751_;
  wire _1752_;
  wire _1753_;
  wire _1754_;
  wire _1755_;
  wire _1756_;
  wire _1757_;
  wire _1758_;
  wire _1759_;
  wire _1760_;
  wire _1761_;
  wire _1762_;
  wire _1763_;
  wire _1764_;
  wire _1765_;
  wire _1766_;
  wire _1767_;
  wire _1768_;
  wire _1769_;
  wire _1770_;
  wire _1771_;
  wire _1772_;
  wire _1773_;
  wire _1774_;
  wire _1775_;
  wire _1776_;
  wire _1777_;
  wire _1778_;
  wire _1779_;
  wire _1780_;
  wire _1781_;
  wire _1782_;
  wire _1783_;
  wire _1784_;
  wire _1785_;
  wire _1786_;
  wire _1787_;
  wire _1788_;
  wire _1789_;
  wire _1790_;
  wire _1791_;
  wire _1792_;
  wire _1793_;
  wire _1794_;
  wire _1795_;
  wire _1796_;
  wire _1797_;
  wire _1798_;
  wire _1799_;
  wire _1800_;
  wire _1801_;
  wire _1802_;
  wire _1803_;
  wire _1804_;
  wire _1805_;
  wire _1806_;
  wire _1807_;
  wire _1808_;
  wire _1809_;
  wire _1810_;
  wire _1811_;
  wire _1812_;
  wire _1813_;
  wire _1814_;
  wire _1815_;
  wire _1816_;
  wire _1817_;
  wire _1818_;
  wire _1819_;
  wire _1820_;
  wire _1821_;
  wire _1822_;
  wire _1823_;
  wire _1824_;
  wire _1825_;
  wire _1826_;
  wire _1827_;
  wire _1828_;
  wire _1829_;
  wire _1830_;
  wire _1831_;
  wire _1832_;
  wire _1833_;
  wire _1834_;
  wire _1835_;
  wire _1836_;
  wire _1837_;
  wire _1838_;
  wire _1839_;
  wire _1840_;
  wire _1841_;
  wire _1842_;
  wire _1843_;
  wire _1844_;
  wire _1845_;
  wire _1846_;
  wire _1847_;
  wire _1848_;
  wire _1849_;
  wire _1850_;
  wire _1851_;
  wire _1852_;
  wire _1853_;
  wire _1854_;
  wire _1855_;
  wire _1856_;
  wire _1857_;
  wire _1858_;
  wire _1859_;
  wire _1860_;
  wire _1861_;
  wire _1862_;
  wire _1863_;
  wire _1864_;
  wire _1865_;
  wire _1866_;
  wire _1867_;
  wire _1868_;
  wire _1869_;
  wire _1870_;
  wire _1871_;
  wire _1872_;
  wire _1873_;
  wire _1874_;
  wire _1875_;
  wire _1876_;
  wire _1877_;
  wire _1878_;
  wire _1879_;
  wire _1880_;
  wire _1881_;
  wire _1882_;
  wire _1883_;
  wire _1884_;
  wire _1885_;
  wire _1886_;
  wire _1887_;
  wire _1888_;
  wire _1889_;
  wire _1890_;
  wire _1891_;
  wire _1892_;
  wire _1893_;
  wire _1894_;
  wire _1895_;
  wire _1896_;
  wire _1897_;
  wire _1898_;
  wire _1899_;
  wire _1900_;
  wire _1901_;
  wire _1902_;
  wire _1903_;
  wire _1904_;
  wire _1905_;
  wire _1906_;
  wire _1907_;
  wire _1908_;
  wire _1909_;
  wire _1910_;
  wire _1911_;
  wire _1912_;
  wire _1913_;
  wire _1914_;
  wire _1915_;
  wire _1916_;
  wire _1917_;
  wire _1918_;
  wire _1919_;
  wire _1920_;
  wire _1921_;
  wire _1922_;
  wire _1923_;
  wire _1924_;
  wire _1925_;
  wire _1926_;
  wire _1927_;
  wire _1928_;
  wire _1929_;
  wire _1930_;
  wire _1931_;
  wire _1932_;
  wire _1933_;
  wire _1934_;
  wire _1935_;
  wire _1936_;
  wire _1937_;
  wire _1938_;
  wire _1939_;
  wire _1940_;
  wire _1941_;
  wire _1942_;
  wire _1943_;
  wire _1944_;
  wire _1945_;
  wire _1946_;
  wire _1947_;
  wire _1948_;
  wire _1949_;
  wire _1950_;
  wire _1951_;
  wire _1952_;
  wire _1953_;
  wire _1954_;
  wire _1955_;
  wire _1956_;
  wire _1957_;
  wire _1958_;
  wire _1959_;
  wire _1960_;
  wire _1961_;
  wire _1962_;
  wire _1963_;
  wire _1964_;
  wire _1965_;
  wire _1966_;
  wire _1967_;
  wire _1968_;
  wire _1969_;
  wire _1970_;
  wire _1971_;
  wire _1972_;
  wire _1973_;
  wire _1974_;
  wire _1975_;
  wire _1976_;
  wire _1977_;
  wire _1978_;
  wire _1979_;
  wire _1980_;
  wire _1981_;
  wire _1982_;
  wire _1983_;
  wire _1984_;
  wire _1985_;
  wire _1986_;
  wire _1987_;
  wire _1988_;
  wire _1989_;
  wire _1990_;
  wire _1991_;
  wire _1992_;
  wire _1993_;
  wire _1994_;
  wire _1995_;
  wire _1996_;
  wire _1997_;
  wire _1998_;
  wire _1999_;
  wire _2000_;
  wire _2001_;
  wire _2002_;
  wire _2003_;
  wire _2004_;
  wire _2005_;
  wire _2006_;
  wire _2007_;
  wire _2008_;
  wire _2009_;
  wire _2010_;
  wire _2011_;
  wire _2012_;
  wire _2013_;
  wire _2014_;
  wire _2015_;
  wire _2016_;
  wire _2017_;
  wire _2018_;
  wire _2019_;
  wire _2020_;
  wire _2021_;
  wire _2022_;
  wire _2023_;
  wire _2024_;
  wire _2025_;
  wire _2026_;
  wire _2027_;
  wire _2028_;
  wire _2029_;
  wire _2030_;
  wire _2031_;
  wire _2032_;
  wire _2033_;
  wire _2034_;
  wire _2035_;
  wire _2036_;
  wire _2037_;
  wire _2038_;
  wire _2039_;
  wire _2040_;
  wire _2041_;
  wire _2042_;
  wire _2043_;
  wire _2044_;
  wire _2045_;
  wire _2046_;
  wire _2047_;
  wire _2048_;
  wire _2049_;
  wire _2050_;
  wire _2051_;
  wire _2052_;
  wire _2053_;
  wire _2054_;
  wire _2055_;
  wire _2056_;
  wire _2057_;
  wire _2058_;
  wire _2059_;
  wire _2060_;
  wire _2061_;
  wire _2062_;
  wire _2063_;
  wire _2064_;
  wire _2065_;
  wire _2066_;
  wire _2067_;
  wire _2068_;
  wire _2069_;
  wire _2070_;
  wire _2071_;
  wire _2072_;
  wire _2073_;
  wire _2074_;
  wire _2075_;
  wire _2076_;
  wire _2077_;
  wire _2078_;
  wire _2079_;
  wire _2080_;
  wire _2081_;
  wire _2082_;
  wire _2083_;
  wire _2084_;
  wire _2085_;
  wire _2086_;
  wire _2087_;
  wire _2088_;
  wire _2089_;
  wire _2090_;
  wire _2091_;
  wire _2092_;
  wire _2093_;
  wire _2094_;
  wire _2095_;
  wire _2096_;
  wire _2097_;
  wire _2098_;
  wire _2099_;
  wire _2100_;
  wire _2101_;
  wire _2102_;
  wire _2103_;
  wire _2104_;
  wire _2105_;
  wire _2106_;
  wire _2107_;
  wire _2108_;
  wire _2109_;
  wire _2110_;
  wire _2111_;
  wire _2112_;
  wire _2113_;
  wire _2114_;
  wire _2115_;
  wire _2116_;
  wire _2117_;
  wire _2118_;
  wire _2119_;
  wire _2120_;
  wire _2121_;
  wire _2122_;
  wire _2123_;
  wire _2124_;
  wire _2125_;
  wire _2126_;
  wire _2127_;
  wire _2128_;
  wire _2129_;
  wire _2130_;
  wire _2131_;
  wire _2132_;
  wire _2133_;
  wire _2134_;
  wire _2135_;
  wire _2136_;
  wire _2137_;
  wire _2138_;
  wire _2139_;
  wire _2140_;
  wire _2141_;
  wire _2142_;
  wire _2143_;
  wire _2144_;
  wire _2145_;
  wire _2146_;
  wire _2147_;
  wire _2148_;
  wire _2149_;
  wire _2150_;
  wire _2151_;
  wire _2152_;
  wire _2153_;
  wire _2154_;
  wire _2155_;
  wire _2156_;
  wire _2157_;
  wire _2158_;
  wire _2159_;
  wire _2160_;
  wire _2161_;
  wire _2162_;
  wire _2163_;
  wire _2164_;
  wire _2165_;
  wire _2166_;
  wire _2167_;
  wire _2168_;
  wire _2169_;
  wire _2170_;
  wire _2171_;
  wire _2172_;
  wire _2173_;
  wire _2174_;
  wire _2175_;
  wire _2176_;
  wire _2177_;
  wire _2178_;
  wire _2179_;
  wire _2180_;
  wire _2181_;
  wire _2182_;
  wire _2183_;
  wire _2184_;
  wire _2185_;
  wire _2186_;
  wire _2187_;
  wire _2188_;
  wire _2189_;
  wire _2190_;
  wire _2191_;
  wire _2192_;
  wire _2193_;
  wire _2194_;
  wire _2195_;
  wire _2196_;
  wire _2197_;
  wire _2198_;
  wire _2199_;
  wire _2200_;
  wire _2201_;
  wire _2202_;
  wire _2203_;
  wire _2204_;
  wire _2205_;
  wire _2206_;
  wire _2207_;
  wire _2208_;
  wire _2209_;
  wire _2210_;
  wire _2211_;
  wire _2212_;
  wire _2213_;
  wire _2214_;
  wire _2215_;
  wire _2216_;
  wire _2217_;
  wire _2218_;
  wire _2219_;
  wire _2220_;
  wire _2221_;
  wire _2222_;
  wire _2223_;
  wire _2224_;
  wire _2225_;
  wire _2226_;
  wire _2227_;
  wire _2228_;
  wire _2229_;
  wire _2230_;
  wire _2231_;
  wire _2232_;
  wire _2233_;
  wire _2234_;
  wire _2235_;
  wire _2236_;
  wire _2237_;
  wire _2238_;
  wire _2239_;
  wire _2240_;
  wire _2241_;
  wire _2242_;
  wire _2243_;
  wire _2244_;
  wire _2245_;
  wire _2246_;
  wire _2247_;
  wire _2248_;
  wire _2249_;
  wire _2250_;
  wire _2251_;
  wire _2252_;
  wire _2253_;
  wire _2254_;
  wire _2255_;
  wire _2256_;
  wire _2257_;
  wire _2258_;
  wire _2259_;
  wire _2260_;
  wire _2261_;
  wire _2262_;
  wire _2263_;
  wire _2264_;
  wire _2265_;
  wire _2266_;
  wire _2267_;
  wire _2268_;
  wire _2269_;
  wire _2270_;
  wire _2271_;
  wire _2272_;
  wire _2273_;
  wire _2274_;
  wire _2275_;
  wire _2276_;
  wire _2277_;
  wire _2278_;
  wire _2279_;
  wire _2280_;
  wire _2281_;
  wire _2282_;
  wire _2283_;
  wire _2284_;
  wire _2285_;
  wire _2286_;
  wire _2287_;
  wire _2288_;
  wire _2289_;
  wire _2290_;
  wire _2291_;
  wire _2292_;
  wire _2293_;
  wire _2294_;
  wire _2295_;
  wire _2296_;
  wire _2297_;
  wire _2298_;
  wire _2299_;
  wire _2300_;
  wire _2301_;
  wire _2302_;
  wire _2303_;
  wire _2304_;
  wire _2305_;
  wire _2306_;
  wire _2307_;
  wire _2308_;
  wire _2309_;
  wire _2310_;
  wire _2311_;
  wire _2312_;
  wire _2313_;
  wire _2314_;
  wire _2315_;
  wire _2316_;
  wire _2317_;
  wire _2318_;
  wire _2319_;
  wire _2320_;
  wire _2321_;
  wire _2322_;
  wire _2323_;
  wire _2324_;
  wire _2325_;
  wire _2326_;
  wire _2327_;
  wire _2328_;
  wire _2329_;
  wire _2330_;
  wire _2331_;
  wire _2332_;
  wire _2333_;
  wire _2334_;
  wire _2335_;
  wire _2336_;
  wire _2337_;
  wire _2338_;
  wire _2339_;
  wire _2340_;
  wire _2341_;
  wire _2342_;
  wire _2343_;
  wire _2344_;
  wire _2345_;
  wire _2346_;
  wire _2347_;
  wire _2348_;
  wire _2349_;
  wire _2350_;
  wire _2351_;
  wire _2352_;
  wire _2353_;
  wire _2354_;
  wire _2355_;
  wire _2356_;
  wire _2357_;
  wire _2358_;
  wire _2359_;
  wire _2360_;
  wire _2361_;
  wire _2362_;
  wire _2363_;
  wire _2364_;
  wire _2365_;
  wire _2366_;
  wire _2367_;
  wire _2368_;
  wire _2369_;
  wire _2370_;
  wire _2371_;
  wire _2372_;
  wire _2373_;
  wire _2374_;
  wire _2375_;
  wire _2376_;
  wire _2377_;
  wire _2378_;
  wire _2379_;
  wire _2380_;
  wire _2381_;
  wire _2382_;
  wire _2383_;
  wire _2384_;
  wire _2385_;
  wire _2386_;
  wire _2387_;
  wire _2388_;
  wire _2389_;
  wire _2390_;
  wire _2391_;
  wire _2392_;
  wire _2393_;
  wire _2394_;
  wire _2395_;
  wire _2396_;
  wire _2397_;
  wire _2398_;
  wire _2399_;
  wire _2400_;
  wire _2401_;
  wire _2402_;
  wire _2403_;
  wire _2404_;
  wire _2405_;
  wire _2406_;
  wire _2407_;
  wire _2408_;
  wire _2409_;
  wire _2410_;
  wire _2411_;
  wire _2412_;
  wire _2413_;
  wire _2414_;
  wire _2415_;
  wire _2416_;
  wire _2417_;
  wire _2418_;
  wire _2419_;
  wire _2420_;
  wire _2421_;
  wire _2422_;
  wire _2423_;
  wire _2424_;
  wire _2425_;
  wire _2426_;
  wire _2427_;
  wire _2428_;
  wire _2429_;
  wire _2430_;
  wire _2431_;
  wire _2432_;
  wire _2433_;
  wire _2434_;
  wire _2435_;
  wire _2436_;
  wire _2437_;
  wire _2438_;
  wire _2439_;
  wire _2440_;
  wire _2441_;
  wire _2442_;
  wire _2443_;
  wire _2444_;
  wire _2445_;
  wire _2446_;
  wire _2447_;
  wire _2448_;
  wire _2449_;
  wire _2450_;
  wire _2451_;
  wire _2452_;
  wire _2453_;
  wire _2454_;
  wire _2455_;
  wire _2456_;
  wire _2457_;
  wire _2458_;
  wire _2459_;
  wire _2460_;
  wire _2461_;
  wire _2462_;
  wire _2463_;
  wire _2464_;
  wire _2465_;
  wire _2466_;
  wire _2467_;
  wire _2468_;
  wire _2469_;
  wire _2470_;
  wire _2471_;
  wire _2472_;
  wire _2473_;
  wire _2474_;
  wire _2475_;
  wire _2476_;
  wire _2477_;
  wire _2478_;
  wire _2479_;
  wire _2480_;
  wire _2481_;
  wire _2482_;
  wire _2483_;
  wire _2484_;
  wire _2485_;
  wire _2486_;
  wire _2487_;
  wire _2488_;
  wire _2489_;
  wire _2490_;
  wire _2491_;
  wire _2492_;
  wire _2493_;
  wire _2494_;
  wire _2495_;
  wire _2496_;
  wire _2497_;
  wire _2498_;
  wire _2499_;
  wire _2500_;
  wire _2501_;
  wire _2502_;
  wire _2503_;
  wire _2504_;
  wire _2505_;
  wire _2506_;
  wire _2507_;
  wire _2508_;
  wire _2509_;
  wire _2510_;
  wire _2511_;
  wire _2512_;
  wire _2513_;
  wire _2514_;
  wire _2515_;
  wire _2516_;
  wire _2517_;
  wire _2518_;
  wire _2519_;
  wire _2520_;
  wire _2521_;
  wire _2522_;
  wire _2523_;
  wire _2524_;
  wire _2525_;
  wire _2526_;
  wire _2527_;
  wire _2528_;
  wire _2529_;
  wire _2530_;
  wire _2531_;
  wire _2532_;
  wire _2533_;
  wire _2534_;
  wire _2535_;
  wire _2536_;
  wire _2537_;
  wire _2538_;
  wire _2539_;
  wire _2540_;
  wire _2541_;
  wire _2542_;
  wire _2543_;
  wire _2544_;
  wire _2545_;
  wire _2546_;
  wire _2547_;
  wire _2548_;
  wire _2549_;
  wire _2550_;
  wire _2551_;
  wire _2552_;
  wire _2553_;
  wire _2554_;
  wire _2555_;
  wire _2556_;
  wire _2557_;
  wire _2558_;
  wire _2559_;
  wire _2560_;
  wire _2561_;
  wire _2562_;
  wire _2563_;
  wire _2564_;
  wire _2565_;
  wire _2566_;
  wire _2567_;
  wire _2568_;
  wire _2569_;
  wire _2570_;
  wire _2571_;
  wire _2572_;
  wire _2573_;
  wire _2574_;
  wire _2575_;
  wire _2576_;
  wire _2577_;
  wire _2578_;
  wire _2579_;
  wire _2580_;
  wire _2581_;
  wire _2582_;
  wire _2583_;
  wire _2584_;
  wire _2585_;
  wire _2586_;
  wire _2587_;
  wire _2588_;
  wire _2589_;
  wire _2590_;
  wire _2591_;
  wire _2592_;
  wire _2593_;
  wire _2594_;
  wire _2595_;
  wire _2596_;
  wire _2597_;
  wire _2598_;
  wire _2599_;
  wire _2600_;
  wire _2601_;
  wire _2602_;
  wire _2603_;
  wire _2604_;
  wire _2605_;
  wire _2606_;
  wire _2607_;
  wire _2608_;
  wire _2609_;
  wire _2610_;
  wire _2611_;
  wire _2612_;
  wire _2613_;
  wire _2614_;
  wire _2615_;
  wire _2616_;
  wire _2617_;
  wire _2618_;
  wire _2619_;
  wire _2620_;
  wire _2621_;
  wire _2622_;
  wire _2623_;
  wire _2624_;
  wire _2625_;
  wire _2626_;
  wire _2627_;
  wire _2628_;
  wire _2629_;
  wire _2630_;
  wire _2631_;
  wire _2632_;
  wire _2633_;
  wire _2634_;
  wire _2635_;
  wire _2636_;
  wire _2637_;
  wire _2638_;
  wire _2639_;
  wire _2640_;
  wire _2641_;
  wire _2642_;
  wire _2643_;
  wire _2644_;
  wire _2645_;
  wire _2646_;
  wire _2647_;
  wire _2648_;
  wire _2649_;
  wire _2650_;
  wire _2651_;
  wire _2652_;
  wire _2653_;
  wire _2654_;
  wire _2655_;
  wire _2656_;
  wire _2657_;
  wire _2658_;
  wire _2659_;
  wire _2660_;
  wire _2661_;
  wire _2662_;
  wire _2663_;
  wire _2664_;
  wire _2665_;
  wire _2666_;
  wire _2667_;
  wire _2668_;
  wire _2669_;
  wire _2670_;
  wire _2671_;
  wire _2672_;
  wire _2673_;
  wire _2674_;
  wire _2675_;
  wire _2676_;
  wire _2677_;
  wire _2678_;
  wire _2679_;
  wire _2680_;
  wire _2681_;
  wire _2682_;
  wire _2683_;
  wire _2684_;
  wire _2685_;
  wire _2686_;
  wire _2687_;
  wire _2688_;
  wire _2689_;
  wire _2690_;
  wire _2691_;
  wire _2692_;
  wire _2693_;
  wire _2694_;
  wire _2695_;
  wire _2696_;
  wire _2697_;
  wire _2698_;
  wire _2699_;
  wire _2700_;
  wire _2701_;
  wire _2702_;
  wire _2703_;
  wire _2704_;
  wire _2705_;
  wire _2706_;
  wire _2707_;
  wire _2708_;
  wire _2709_;
  wire _2710_;
  wire _2711_;
  wire _2712_;
  wire _2713_;
  wire _2714_;
  wire _2715_;
  wire _2716_;
  wire _2717_;
  wire _2718_;
  wire _2719_;
  wire _2720_;
  wire _2721_;
  wire _2722_;
  wire _2723_;
  wire _2724_;
  wire _2725_;
  wire _2726_;
  wire _2727_;
  wire _2728_;
  wire _2729_;
  wire _2730_;
  wire _2731_;
  wire _2732_;
  wire _2733_;
  wire _2734_;
  wire _2735_;
  wire _2736_;
  wire _2737_;
  wire _2738_;
  wire _2739_;
  wire _2740_;
  wire _2741_;
  wire _2742_;
  wire _2743_;
  wire _2744_;
  wire _2745_;
  wire _2746_;
  wire _2747_;
  wire _2748_;
  wire _2749_;
  wire _2750_;
  wire _2751_;
  wire _2752_;
  wire _2753_;
  wire _2754_;
  wire _2755_;
  wire _2756_;
  wire _2757_;
  wire _2758_;
  wire _2759_;
  wire _2760_;
  wire _2761_;
  wire _2762_;
  wire _2763_;
  wire _2764_;
  wire _2765_;
  wire _2766_;
  wire _2767_;
  wire _2768_;
  wire _2769_;
  wire _2770_;
  wire _2771_;
  wire _2772_;
  wire _2773_;
  wire _2774_;
  wire _2775_;
  wire _2776_;
  wire _2777_;
  wire _2778_;
  wire _2779_;
  wire _2780_;
  wire _2781_;
  wire _2782_;
  wire _2783_;
  wire _2784_;
  wire _2785_;
  wire _2786_;
  wire _2787_;
  wire _2788_;
  wire _2789_;
  wire _2790_;
  wire _2791_;
  wire _2792_;
  wire _2793_;
  wire _2794_;
  wire _2795_;
  wire _2796_;
  wire _2797_;
  wire _2798_;
  wire _2799_;
  wire _2800_;
  wire _2801_;
  wire _2802_;
  wire _2803_;
  wire _2804_;
  wire _2805_;
  wire _2806_;
  wire _2807_;
  wire _2808_;
  wire _2809_;
  wire _2810_;
  wire _2811_;
  wire _2812_;
  wire _2813_;
  wire _2814_;
  wire _2815_;
  wire _2816_;
  wire _2817_;
  wire _2818_;
  wire _2819_;
  wire _2820_;
  wire _2821_;
  wire _2822_;
  wire _2823_;
  wire _2824_;
  wire _2825_;
  wire _2826_;
  wire _2827_;
  wire _2828_;
  wire _2829_;
  wire _2830_;
  wire _2831_;
  wire _2832_;
  wire _2833_;
  wire _2834_;
  wire _2835_;
  wire _2836_;
  wire _2837_;
  wire _2838_;
  wire _2839_;
  wire _2840_;
  wire _2841_;
  wire _2842_;
  wire _2843_;
  wire _2844_;
  wire _2845_;
  wire _2846_;
  wire _2847_;
  wire _2848_;
  wire _2849_;
  wire _2850_;
  wire _2851_;
  wire _2852_;
  wire _2853_;
  wire _2854_;
  wire _2855_;
  wire _2856_;
  wire _2857_;
  wire _2858_;
  wire _2859_;
  wire _2860_;
  wire _2861_;
  wire _2862_;
  wire _2863_;
  wire _2864_;
  wire _2865_;
  wire _2866_;
  wire _2867_;
  wire _2868_;
  wire _2869_;
  wire _2870_;
  wire _2871_;
  wire _2872_;
  wire _2873_;
  wire _2874_;
  wire _2875_;
  wire _2876_;
  wire _2877_;
  wire _2878_;
  wire _2879_;
  wire _2880_;
  wire _2881_;
  wire _2882_;
  wire _2883_;
  wire _2884_;
  wire _2885_;
  wire _2886_;
  wire _2887_;
  wire _2888_;
  wire _2889_;
  wire _2890_;
  wire _2891_;
  wire _2892_;
  wire _2893_;
  wire _2894_;
  wire _2895_;
  wire _2896_;
  wire _2897_;
  wire _2898_;
  wire _2899_;
  wire _2900_;
  wire _2901_;
  wire _2902_;
  wire _2903_;
  wire _2904_;
  wire _2905_;
  wire _temp0_;
  wire _temp1_;
  wire _temp2_;
  wire _temp3_;
  wire _temp4_;
  wire _temp5_;
  wire _temp6_;
  wire _temp7_;
  wire _temp8_;
  wire _temp9_;
  wire _temp10_;
  wire _temp11_;
  wire _temp12_;
  wire _temp13_;
  wire _temp14_;
  wire _temp15_;
  wire _temp16_;
  wire _temp17_;
  wire _temp18_;
  wire _temp19_;
  wire _temp20_;
  wire _temp21_;
  wire _temp22_;
  wire _temp23_;
  wire _temp24_;
  wire _temp25_;
  wire _temp26_;
  wire _temp27_;
  wire _temp28_;
  wire _temp29_;
  wire _temp30_;
  wire _temp31_;
  wire _temp32_;
  wire _temp33_;
  wire _temp34_;
  wire _temp35_;
  wire _temp36_;
  wire _temp37_;
  wire _temp38_;
  wire _temp39_;
  wire _temp40_;
  wire _temp41_;
  wire _temp42_;
  wire _temp43_;
  wire _temp44_;
  wire _temp45_;
  wire _temp46_;
  wire _temp47_;
  wire _temp48_;
  wire _temp49_;
  wire _temp50_;
  wire _temp51_;
  wire _temp52_;
  wire _temp53_;
  wire _temp54_;
  wire _temp55_;
  wire _temp56_;
  wire _temp57_;
  wire _temp58_;
  wire _temp59_;
  wire _temp60_;
  wire _temp61_;
  wire _temp62_;
  wire _temp63_;
  wire _temp64_;
  wire _temp65_;
  wire _temp66_;
  wire _temp67_;
  wire _temp68_;
  wire _temp69_;
  wire _temp70_;
  wire _temp71_;
  wire _temp72_;
  wire _temp73_;
  wire _temp74_;
  wire _temp75_;
  wire _temp76_;
  wire _temp77_;
  wire _temp78_;
  wire _temp79_;
  wire _temp80_;
  wire _temp81_;
  wire _temp82_;
  wire _temp83_;
  wire _temp84_;
  wire _temp85_;
  wire _temp86_;
  wire _temp87_;
  wire _temp88_;
  wire _temp89_;
  wire _temp90_;
  wire _temp91_;
  wire _temp92_;
  wire _temp93_;
  wire _temp94_;
  wire _temp95_;
  wire _temp96_;
  wire _temp97_;
  wire _temp98_;
  wire _temp99_;
  wire _temp100_;
  wire _temp101_;
  wire _temp102_;
  wire _temp103_;
  wire _temp104_;
  wire _temp105_;
  wire _temp106_;
  wire _temp107_;
  wire _temp108_;
  wire _temp109_;
  wire _temp110_;
  wire _temp111_;
  wire _temp112_;
  wire _temp113_;
  wire _temp114_;
  wire _temp115_;
  wire _temp116_;
  wire _temp117_;
  wire _temp118_;
  wire _temp119_;
  wire _temp120_;
  wire _temp121_;
  wire _temp122_;
  wire _temp123_;
  wire _temp124_;
  wire _temp125_;
  wire _temp126_;
  wire _temp127_;
  wire _temp128_;
  wire _temp129_;
  wire _temp130_;
  wire _temp131_;
  wire _temp132_;
  wire _temp133_;
  wire _temp134_;
  wire _temp135_;
  wire _temp136_;
  wire _temp137_;
  wire _temp138_;
  wire _temp139_;
  wire _temp140_;
  wire _temp141_;
  wire _temp142_;
  wire _temp143_;
  wire _temp144_;
  wire _temp145_;
  wire _temp146_;
  wire _temp147_;
  wire _temp148_;
  wire _temp149_;
  wire _temp150_;
  wire _temp151_;
  wire _temp152_;
  wire _temp153_;
  wire _temp154_;
  wire _temp155_;
  wire _temp156_;
  wire _temp157_;
  wire _temp158_;
  wire _temp159_;
  wire _temp160_;
  wire _temp161_;
  wire _temp162_;
  wire _temp163_;
  wire _temp164_;
  wire _temp165_;
  wire _temp166_;
  wire _temp167_;
  wire _temp168_;
  wire _temp169_;
  wire _temp170_;
  wire _temp171_;
  wire _temp172_;
  wire _temp173_;
  wire _temp174_;
  wire _temp175_;
  wire _temp176_;
  wire _temp177_;
  wire _temp178_;
  wire _temp179_;
  wire _temp180_;
  wire _temp181_;
  wire _temp182_;
  wire _temp183_;
  wire _temp184_;
  wire _temp185_;
  wire _temp186_;
  wire _temp187_;
  wire _temp188_;
  wire _temp189_;
  wire _temp190_;
  wire _temp191_;
  wire _temp192_;
  wire _temp193_;
  wire _temp194_;
  wire _temp195_;
  wire _temp196_;
  wire _temp197_;
  wire _temp198_;
  wire _temp199_;
  wire _temp200_;
  wire _temp201_;
  wire _temp202_;
  wire _temp203_;
  wire _temp204_;
  wire _temp205_;
  wire _temp206_;
  wire _temp207_;
  wire _temp208_;
  wire _temp209_;
  wire _temp210_;
  wire _temp211_;
  wire _temp212_;
  wire _temp213_;
  wire _temp214_;
  wire _temp215_;
  wire _temp216_;
  wire _temp217_;
  wire _temp218_;
  wire _temp219_;
  wire _temp220_;
  wire _temp221_;
  wire _temp222_;
  wire _temp223_;
  wire _temp224_;
  wire _temp225_;
  wire _temp226_;
  wire _temp227_;
  wire _temp228_;
  wire _temp229_;
  wire _temp230_;
  wire _temp231_;
  wire _temp232_;
  wire _temp233_;
  wire _temp234_;
  wire _temp235_;
  wire _temp236_;
  wire _temp237_;
  wire _temp238_;
  wire _temp239_;
  wire _temp240_;
  wire _temp241_;
  wire _temp242_;
  wire _temp243_;
  wire _temp244_;
  wire _temp245_;
  wire _temp246_;
  wire _temp247_;
  wire _temp248_;
  wire _temp249_;
  wire _temp250_;
  wire _temp251_;
  wire _temp252_;
  wire _temp253_;
  wire _temp254_;
  wire _temp255_;
  wire _temp256_;
  wire _temp257_;
  wire _temp258_;
  wire _temp259_;
  wire _temp260_;
  wire _temp261_;
  wire _temp262_;
  wire _temp263_;
  wire _temp264_;
  wire _temp265_;
  wire _temp266_;
  wire _temp267_;
  wire _temp268_;
  wire _temp269_;
  wire _temp270_;
  wire _temp271_;
  wire _temp272_;
  wire _temp273_;
  wire _temp274_;
  wire _temp275_;
  wire _temp276_;
  wire _temp277_;
  wire _temp278_;
  wire _temp279_;
  wire _temp280_;
  wire _temp281_;
  wire _temp282_;
  wire _temp283_;
  wire _temp284_;
  wire _temp285_;
  wire _temp286_;
  wire _temp287_;
  wire _temp288_;
  wire _temp289_;
  wire _temp290_;
  wire _temp291_;
  wire _temp292_;
  wire _temp293_;
  wire _temp294_;
  wire _temp295_;
  wire _temp296_;
  wire _temp297_;
  wire _temp298_;
  wire _temp299_;
  wire _temp300_;
  wire _temp301_;
  wire _temp302_;
  wire _temp303_;
  wire _temp304_;
  wire _temp305_;
  wire _temp306_;
  wire _temp307_;
  wire _temp308_;
  wire _temp309_;
  wire _temp310_;
  wire _temp311_;
  wire _temp312_;
  wire _temp313_;
  wire _temp314_;
  wire _temp315_;
  wire _temp316_;
  wire _temp317_;
  wire _temp318_;
  wire _temp319_;
  wire _temp320_;
  wire _temp321_;
  wire _temp322_;
  wire _temp323_;
  wire _temp324_;
  wire _temp325_;
  wire _temp326_;
  wire _temp327_;
  wire _temp328_;
  wire _temp329_;
  wire _temp330_;
  wire _temp331_;
  wire _temp332_;
  wire _temp333_;
  wire _temp334_;
  wire _temp335_;
  wire _temp336_;
  wire _temp337_;
  wire _temp338_;
  wire _temp339_;
  wire _temp340_;
  wire _temp341_;
  wire _temp342_;
  wire _temp343_;
  wire _temp344_;
  wire _temp345_;
  wire _temp346_;
  wire _temp347_;
  wire _temp348_;
  wire _temp349_;
  wire _temp350_;
  wire _temp351_;
  wire _temp352_;
  wire _temp353_;
  wire _temp354_;
  wire _temp355_;
  wire _temp356_;
  wire _temp357_;
  wire _temp358_;
  wire _temp359_;
  wire _temp360_;
  wire _temp361_;
  wire _temp362_;
  wire _temp363_;
  wire _temp364_;
  wire _temp365_;
  wire _temp366_;
  wire _temp367_;
  wire _temp368_;
  wire _temp369_;
  wire _temp370_;
  wire _temp371_;
  wire _temp372_;
  wire _temp373_;
  wire _temp374_;
  wire _temp375_;
  wire _temp376_;
  wire _temp377_;
  wire _temp378_;
  wire _temp379_;
  wire _temp380_;
  wire _temp381_;
  wire _temp382_;
  wire _temp383_;
  wire _temp384_;
  wire _temp385_;
  wire _temp386_;
  wire _temp387_;
  wire _temp388_;
  wire _temp389_;
  wire _temp390_;
  wire _temp391_;
  wire _temp392_;
  wire _temp393_;
  wire _temp394_;
  wire _temp395_;
  wire _temp396_;
  wire _temp397_;
  wire _temp398_;
  wire _temp399_;
  wire _temp400_;
  wire _temp401_;
  wire _temp402_;
  wire _temp403_;
  wire _temp404_;
  wire _temp405_;
  wire _temp406_;
  wire _temp407_;
  wire _temp408_;
  wire _temp409_;
  wire _temp410_;
  wire _temp411_;
  wire _temp412_;
  wire _temp413_;
  wire _temp414_;
  wire _temp415_;
  wire _temp416_;
  wire _temp417_;
  wire _temp418_;
  wire _temp419_;
  wire _temp420_;
  wire _temp421_;
  wire _temp422_;
  wire _temp423_;
  wire _temp424_;
  wire _temp425_;
  wire _temp426_;
  wire _temp427_;
  wire _temp428_;
  wire _temp429_;
  wire _temp430_;
  wire _temp431_;
  wire _temp432_;
  wire _temp433_;
  wire _temp434_;
  wire _temp435_;
  wire _temp436_;
  wire _temp437_;
  wire _temp438_;
  wire _temp439_;
  wire _temp440_;
  wire _temp441_;
  wire _temp442_;
  wire _temp443_;
  wire _temp444_;
  wire _temp445_;
  wire _temp446_;
  wire _temp447_;
  wire _temp448_;
  wire _temp449_;
  wire _temp450_;
  wire _temp451_;
  wire _temp452_;
  wire _temp453_;
  wire _temp454_;
  wire _temp455_;
  wire _temp456_;
  wire _temp457_;
  wire _temp458_;
  wire _temp459_;
  wire _temp460_;
  wire _temp461_;
  wire _temp462_;
  wire _temp463_;
  wire _temp464_;
  wire _temp465_;
  wire _temp466_;
  wire _temp467_;
  wire _temp468_;
  wire _temp469_;
  wire _temp470_;
  wire _temp471_;
  wire _temp472_;
  wire _temp473_;
  wire _temp474_;
  wire _temp475_;
  wire _temp476_;
  wire _temp477_;
  wire _temp478_;
  wire _temp479_;
  wire _temp480_;
  wire _temp481_;
  wire _temp482_;
  wire _temp483_;
  wire _temp484_;
  wire _temp485_;
  wire _temp486_;
  wire _temp487_;
  wire _temp488_;
  wire _temp489_;
  wire _temp490_;
  wire _temp491_;
  wire _temp492_;
  wire _temp493_;
  wire _temp494_;
  wire _temp495_;
  wire _temp496_;
  wire _temp497_;
  wire _temp498_;
  wire _temp499_;
  wire _temp500_;
  wire _temp501_;
  wire _temp502_;
  wire _temp503_;
  wire _temp504_;
  wire _temp505_;
  wire _temp506_;
  wire _temp507_;
  wire _temp508_;
  wire _temp509_;
  wire _temp510_;
  wire _temp511_;
  wire _temp512_;
  wire _temp513_;
  wire _temp514_;
  wire _temp515_;
  wire _temp516_;
  wire _temp517_;
  wire _temp518_;
  wire _temp519_;
  wire _temp520_;
  wire _temp521_;
  wire _temp522_;
  wire _temp523_;
  wire _temp524_;
  wire _temp525_;
  wire _temp526_;
  wire _temp527_;
  wire _temp528_;
  wire _temp529_;
  wire _temp530_;
  wire _temp531_;
  wire _temp532_;
  wire _temp533_;
  wire _temp534_;
  wire _temp535_;
  wire _temp536_;
  wire _temp537_;
  wire _temp538_;
  wire _temp539_;
  wire _temp540_;
  wire _temp541_;
  wire _temp542_;
  wire _temp543_;
  wire _temp544_;
  wire _temp545_;
  wire _temp546_;
  wire _temp547_;
  wire _temp548_;
  wire _temp549_;
  wire _temp550_;
  wire _temp551_;
  wire _temp552_;
  wire _temp553_;
  wire _temp554_;
  wire _temp555_;
  wire _temp556_;
  wire _temp557_;
  wire _temp558_;
  wire _temp559_;
  wire _temp560_;
  wire _temp561_;
  wire _temp562_;
  wire _temp563_;
  wire _temp564_;
  wire _temp565_;
  wire _temp566_;
  wire _temp567_;
  wire _temp568_;
  wire _temp569_;
  wire _temp570_;
  wire _temp571_;
  wire _temp572_;
  wire _temp573_;
  wire _temp574_;
  wire _temp575_;
  wire _temp576_;
  wire _temp577_;
  wire _temp578_;
  wire _temp579_;
  wire _temp580_;
  wire _temp581_;
  wire _temp582_;
  wire _temp583_;
  wire _temp584_;
  wire _temp585_;
  wire _temp586_;
  wire _temp587_;
  wire _temp588_;
  wire _temp589_;
  wire _temp590_;
  wire _temp591_;
  wire _temp592_;
  wire _temp593_;
  wire _temp594_;
  wire _temp595_;
  wire _temp596_;
  wire _temp597_;
  wire _temp598_;
  wire _temp599_;
  wire _temp600_;
  wire _temp601_;
  wire _temp602_;
  wire _temp603_;
  wire _temp604_;
  wire _temp605_;
  wire _temp606_;
  wire _temp607_;
  wire _temp608_;
  wire _temp609_;
  wire _temp610_;
  wire _temp611_;
  wire _temp612_;
  wire _temp613_;
  wire _temp614_;
  wire _temp615_;
  wire _temp616_;
  wire _temp617_;
  wire _temp618_;
  wire _temp619_;
  wire _temp620_;
  wire _temp621_;
  wire _temp622_;
  wire _temp623_;
  wire _temp624_;
  wire _temp625_;
  wire _temp626_;
  wire _temp627_;
  wire _temp628_;
  wire _temp629_;
  wire _temp630_;
  wire _temp631_;
  wire _temp632_;
  wire _temp633_;
  wire _temp634_;
  wire _temp635_;
  wire _temp636_;
  wire _temp637_;
  wire _temp638_;
  wire _temp639_;
  wire _temp640_;
  wire _temp641_;
  wire _temp642_;
  wire _temp643_;
  wire _temp644_;
  wire _temp645_;
  wire _temp646_;
  wire _temp647_;
  wire _temp648_;
  wire _temp649_;
  wire _temp650_;
  wire _temp651_;
  wire _temp652_;
  wire _temp653_;
  wire _temp654_;
  wire _temp655_;
  wire _temp656_;
  wire _temp657_;
  wire _temp658_;
  wire _temp659_;
  wire _temp660_;
  wire _temp661_;
  wire _temp662_;
  wire _temp663_;
  wire _temp664_;
  wire _temp665_;
  wire _temp666_;
  wire _temp667_;
  wire _temp668_;
  wire _temp669_;
  wire _temp670_;
  wire _temp671_;
  wire _temp672_;
  wire _temp673_;
  wire _temp674_;
  wire _temp675_;
  wire _temp676_;
  wire _temp677_;
  wire _temp678_;
  wire _temp679_;
  wire _temp680_;
  wire _temp681_;
  wire _temp682_;
  wire _temp683_;
  wire _temp684_;
  wire _temp685_;
  wire _temp686_;
  wire _temp687_;
  wire _temp688_;
  wire _temp689_;
  wire _temp690_;
  wire _temp691_;
  wire _temp692_;
  wire _temp693_;
  wire _temp694_;
  wire _temp695_;
  wire _temp696_;
  wire _temp697_;
  wire _temp698_;
  wire _temp699_;
  wire _temp700_;
  wire _temp701_;
  wire _temp702_;
  wire _temp703_;
  wire _temp704_;
  wire _temp705_;
  wire _temp706_;
  wire _temp707_;
  wire _temp708_;
  wire _temp709_;
  wire _temp710_;
  wire _temp711_;
  wire _temp712_;
  wire _temp713_;
  wire _temp714_;
  wire _temp715_;
  wire _temp716_;
  wire _temp717_;
  wire _temp718_;
  wire _temp719_;
  wire _temp720_;
  wire _temp721_;
  wire _temp722_;
  wire _temp723_;
  wire _temp724_;
  wire _temp725_;
  wire _temp726_;
  wire _temp727_;
  wire _temp728_;
  wire _temp729_;
  wire _temp730_;
  wire _temp731_;
  wire _temp732_;
  wire _temp733_;
  wire _temp734_;
  wire _temp735_;
  wire _temp736_;
  wire _temp737_;
  wire _temp738_;
  wire _temp739_;
  wire _temp740_;
  wire _temp741_;
  wire _temp742_;
  wire _temp743_;
  wire _temp744_;
  wire _temp745_;
  wire _temp746_;
  wire _temp747_;
  wire _temp748_;
  wire _temp749_;
  wire _temp750_;
  wire _temp751_;
  wire _temp752_;
  wire _temp753_;
  wire _temp754_;
  wire _temp755_;
  wire _temp756_;
  wire _temp757_;
  wire _temp758_;
  wire _temp759_;
  wire _temp760_;
  wire _temp761_;
  wire _temp762_;
  wire _temp763_;
  wire _temp764_;
  wire _temp765_;
  wire _temp766_;
  wire _temp767_;
  wire _temp768_;
  wire _temp769_;
  wire _temp770_;
  wire _temp771_;
  wire _temp772_;
  wire _temp773_;
  wire _temp774_;
  wire _temp775_;
  wire _temp776_;
  wire _temp777_;
  wire _temp778_;
  wire _temp779_;
  wire _temp780_;
  wire _temp781_;
  wire _temp782_;
  wire _temp783_;
  wire _temp784_;
  wire _temp785_;
  wire _temp786_;
  wire _temp787_;
  wire _temp788_;
  wire _temp789_;
  wire _temp790_;
  wire _temp791_;
  wire _temp792_;
  wire _temp793_;
  wire _temp794_;
  wire _temp795_;
  wire _temp796_;
  wire _temp797_;
  wire _temp798_;
  wire _temp799_;
  wire _temp800_;
  wire _temp801_;
  wire _temp802_;
  wire _temp803_;
  wire _temp804_;
  wire _temp805_;
  wire _temp806_;
  wire _temp807_;
  wire _temp808_;
  wire _temp809_;
  wire _temp810_;
  wire _temp811_;
  wire _temp812_;
  wire _temp813_;
  wire _temp814_;
  wire _temp815_;
  wire _temp816_;
  wire _temp817_;
  wire _temp818_;
  wire _temp819_;
  wire _temp820_;
  wire _temp821_;
  wire _temp822_;
  wire _temp823_;
  wire _temp824_;
  wire _temp825_;
  wire _temp826_;
  wire _temp827_;
  wire _temp828_;
  wire _temp829_;
  wire _temp830_;
  wire _temp831_;
  wire _temp832_;
  wire _temp833_;
  wire _temp834_;
  wire _temp835_;
  wire _temp836_;
  wire _temp837_;
  wire _temp838_;
  wire _temp839_;
  wire _temp840_;
  wire _temp841_;
  wire _temp842_;
  wire _temp843_;
  wire _temp844_;
  wire _temp845_;
  wire _temp846_;
  wire _temp847_;
  wire _temp848_;
  wire _temp849_;
  wire _temp850_;
  wire _temp851_;
  wire _temp852_;
  wire _temp853_;
  wire _temp854_;
  wire _temp855_;
  wire _temp856_;
  wire _temp857_;
  wire _temp858_;
  wire _temp859_;
  wire _temp860_;
  wire _temp861_;
  wire _temp862_;
  wire _temp863_;
  wire _temp864_;
  wire _temp865_;
  wire _temp866_;
  wire _temp867_;
  wire _temp868_;
  wire _temp869_;
  wire _temp870_;
  wire _temp871_;
  wire _temp872_;
  wire _temp873_;
  wire _temp874_;
  wire _temp875_;
  wire _temp876_;
  wire _temp877_;
  wire _temp878_;
  wire _temp879_;
  wire _temp880_;
  wire _temp881_;
  wire _temp882_;
  wire _temp883_;
  wire _temp884_;
  wire _temp885_;
  wire _temp886_;
  wire _temp887_;
  wire _temp888_;
  wire _temp889_;
  wire _temp890_;
  wire _temp891_;
  wire _temp892_;
  wire _temp893_;
  wire _temp894_;
  wire _temp895_;
  wire _temp896_;
  wire _temp897_;
  wire _temp898_;
  wire _temp899_;
  wire _temp900_;
  wire _temp901_;
  wire _temp902_;
  wire _temp903_;
  wire _temp904_;
  wire _temp905_;
  wire _temp906_;
  wire _temp907_;
  wire _temp908_;
  wire _temp909_;
  wire _temp910_;
  wire _temp911_;
  wire _temp912_;
  wire _temp913_;
  wire _temp914_;
  wire _temp915_;
  wire _temp916_;
  wire _temp917_;
  wire _temp918_;
  wire _temp919_;
  wire _temp920_;
  wire _temp921_;
  wire _temp922_;
  wire _temp923_;
  wire _temp924_;
  wire _temp925_;
  wire _temp926_;
  wire _temp927_;
  wire _temp928_;
  wire _temp929_;
  wire _temp930_;
  wire _temp931_;
  wire _temp932_;
  wire _temp933_;
  wire _temp934_;
  wire _temp935_;
  wire _temp936_;
  wire _temp937_;
  wire _temp938_;
  wire _temp939_;
  wire _temp940_;
  wire _temp941_;
  wire _temp942_;
  wire _temp943_;
  wire _temp944_;
  wire _temp945_;
  wire _temp946_;
  wire _temp947_;
  wire _temp948_;
  wire _temp949_;
  wire _temp950_;
  wire _temp951_;
  wire _temp952_;
  wire _temp953_;
  wire _temp954_;
  wire _temp955_;
  wire _temp956_;
  wire _temp957_;
  wire _temp958_;
  wire _temp959_;
  wire _temp960_;
  wire _temp961_;
  wire _temp962_;
  wire _temp963_;
  wire _temp964_;
  wire _temp965_;
  wire _temp966_;
  wire _temp967_;
  wire _temp968_;
  wire _temp969_;
  wire _temp970_;
  wire _temp971_;
  wire _temp972_;
  wire _temp973_;
  wire _temp974_;
  wire _temp975_;
  wire _temp976_;
  wire _temp977_;
  wire _temp978_;
  wire _temp979_;
  wire _temp980_;
  wire _temp981_;
  wire _temp982_;
  wire _temp983_;
  wire _temp984_;
  wire _temp985_;
  wire _temp986_;
  wire _temp987_;
  wire _temp988_;
  wire _temp989_;
  wire _temp990_;
  wire _temp991_;
  wire _temp992_;
  wire _temp993_;
  wire _temp994_;
  wire _temp995_;
  wire _temp996_;
  wire _temp997_;
  wire _temp998_;
  wire _temp999_;
  wire _temp1000_;
  wire _temp1001_;
  wire _temp1002_;
  wire _temp1003_;
  wire _temp1004_;
  wire _temp1005_;
  wire _temp1006_;
  wire _temp1007_;
  wire _temp1008_;
  wire _temp1009_;
  wire _temp1010_;
  wire _temp1011_;
  wire _temp1012_;
  wire _temp1013_;
  wire _temp1014_;
  wire _temp1015_;
  wire _temp1016_;
  wire _temp1017_;
  wire _temp1018_;
  wire _temp1019_;
  wire _temp1020_;
  wire _temp1021_;
  wire _temp1022_;
  wire _temp1023_;
  wire _temp1024_;
  wire _temp1025_;
  wire _temp1026_;
  wire _temp1027_;
  wire _temp1028_;
  wire _temp1029_;
  wire _temp1030_;
  wire _temp1031_;
  wire _temp1032_;
  wire _temp1033_;
  wire _temp1034_;
  wire _temp1035_;
  wire _temp1036_;
  wire _temp1037_;
  wire _temp1038_;
  wire _temp1039_;
  wire _temp1040_;
  wire _temp1041_;
  wire _temp1042_;
  wire _temp1043_;
  wire _temp1044_;
  wire _temp1045_;
  wire _temp1046_;
  wire _temp1047_;
  wire _temp1048_;
  wire _temp1049_;
  wire _temp1050_;
  wire _temp1051_;
  wire _temp1052_;
  wire _temp1053_;
  wire _temp1054_;
  wire _temp1055_;
  wire _temp1056_;
  wire _temp1057_;
  wire _temp1058_;
  wire _temp1059_;
  wire _temp1060_;
  wire _temp1061_;
  wire _temp1062_;
  wire _temp1063_;
  wire _temp1064_;
  wire _temp1065_;
  wire _temp1066_;
  wire _temp1067_;
  wire _temp1068_;
  wire _temp1069_;
  wire _temp1070_;
  wire _temp1071_;
  wire _temp1072_;
  wire _temp1073_;
  wire _temp1074_;
  wire _temp1075_;
  wire _temp1076_;
  wire _temp1077_;
  wire _temp1078_;
  wire _temp1079_;
  wire _temp1080_;
  wire _temp1081_;
  wire _temp1082_;
  wire _temp1083_;
  wire _temp1084_;
  wire _temp1085_;
  wire _temp1086_;
  wire _temp1087_;
  wire _temp1088_;
  wire _temp1089_;
  wire _temp1090_;
  wire _temp1091_;
  wire _temp1092_;
  wire _temp1093_;
  wire _temp1094_;
  wire _temp1095_;
  wire _temp1096_;
  wire _temp1097_;
  wire _temp1098_;
  wire _temp1099_;
  wire _temp1100_;
  wire _temp1101_;
  wire _temp1102_;
  wire _temp1103_;
  wire _temp1104_;
  wire _temp1105_;
  wire _temp1106_;
  wire _temp1107_;
  wire _temp1108_;
  wire _temp1109_;
  wire _temp1110_;
  wire _temp1111_;
  wire _temp1112_;
  wire _temp1113_;
  wire _temp1114_;
  wire _temp1115_;
  wire _temp1116_;
  wire _temp1117_;
  wire _temp1118_;
  wire _temp1119_;
  wire _temp1120_;
  wire _temp1121_;
  wire _temp1122_;
  wire _temp1123_;
  wire _temp1124_;
  wire _temp1125_;
  wire _temp1126_;
  wire _temp1127_;
  wire _temp1128_;
  wire _temp1129_;
  wire _temp1130_;
  wire _temp1131_;
  wire _temp1132_;
  wire _temp1133_;
  wire _temp1134_;
  wire _temp1135_;
  wire _temp1136_;
  wire _temp1137_;
  wire _temp1138_;
  wire _temp1139_;
  wire _temp1140_;
  wire _temp1141_;
  wire _temp1142_;
  wire _temp1143_;
  wire _temp1144_;
  wire _temp1145_;
  wire _temp1146_;
  wire _temp1147_;
  wire _temp1148_;
  wire _temp1149_;
  wire _temp1150_;
  wire _temp1151_;
  wire _temp1152_;
  wire _temp1153_;
  wire _temp1154_;
  wire _temp1155_;
  wire _temp1156_;
  wire _temp1157_;
  wire _temp1158_;
  wire _temp1159_;
  wire _temp1160_;
  wire _temp1161_;
  wire _temp1162_;
  wire _temp1163_;
  wire _temp1164_;
  wire _temp1165_;
  wire _temp1166_;
  wire _temp1167_;
  wire _temp1168_;
  wire _temp1169_;
  wire _temp1170_;
  wire _temp1171_;
  wire _temp1172_;
  wire _temp1173_;
  wire _temp1174_;
  wire _temp1175_;
  wire _temp1176_;
  wire _temp1177_;
  wire _temp1178_;
  wire _temp1179_;
  wire _temp1180_;
  wire _temp1181_;
  wire _temp1182_;
  wire _temp1183_;
  wire _temp1184_;
  wire _temp1185_;
  wire _temp1186_;
  wire _temp1187_;
  wire _temp1188_;
  wire _temp1189_;
  wire _temp1190_;
  wire _temp1191_;
  wire _temp1192_;
  wire _temp1193_;
  wire _temp1194_;
  wire _temp1195_;
  wire _temp1196_;
  wire _temp1197_;
  wire _temp1198_;
  wire _temp1199_;
  wire _temp1200_;
  wire _temp1201_;
  wire _temp1202_;
  wire _temp1203_;
  wire _temp1204_;
  wire _temp1205_;
  wire _temp1206_;
  wire _temp1207_;
  wire _temp1208_;
  wire _temp1209_;
  wire _temp1210_;
  wire _temp1211_;
  wire _temp1212_;
  wire _temp1213_;
  wire _temp1214_;
  wire _temp1215_;
  wire _temp1216_;
  wire _temp1217_;
  wire _temp1218_;
  wire _temp1219_;
  wire _temp1220_;
  wire _temp1221_;
  wire _temp1222_;
  wire _temp1223_;
  wire _temp1224_;
  wire _temp1225_;
  wire _temp1226_;
  wire _temp1227_;
  wire _temp1228_;
  wire _temp1229_;
  wire _temp1230_;
  wire _temp1231_;
  wire _temp1232_;
  wire _temp1233_;
  wire _temp1234_;
  wire _temp1235_;
  wire _temp1236_;
  wire _temp1237_;
  wire _temp1238_;
  wire _temp1239_;
  wire _temp1240_;
  wire _temp1241_;
  wire _temp1242_;
  wire _temp1243_;
  wire _temp1244_;
  wire _temp1245_;
  wire _temp1246_;
  wire _temp1247_;
  wire _temp1248_;
  wire _temp1249_;
  wire _temp1250_;
  wire _temp1251_;
  wire _temp1252_;
  wire _temp1253_;
  wire _temp1254_;
  wire _temp1255_;
  wire _temp1256_;
  wire _temp1257_;
  wire _temp1258_;
  wire _temp1259_;
  wire _temp1260_;
  wire _temp1261_;
  wire _temp1262_;
  wire _temp1263_;
  wire _temp1264_;
  wire _temp1265_;
  wire _temp1266_;
  wire _temp1267_;
  wire _temp1268_;
  wire _temp1269_;
  wire _temp1270_;
  wire _temp1271_;
  wire _temp1272_;
  wire _temp1273_;
  wire _temp1274_;
  wire _temp1275_;
  wire _temp1276_;
  wire _temp1277_;
  wire _temp1278_;
  wire _temp1279_;
  wire _temp1280_;
  wire _temp1281_;
  wire _temp1282_;
  wire _temp1283_;
  wire _temp1284_;
  wire _temp1285_;
  wire _temp1286_;
  wire _temp1287_;
  wire _temp1288_;
  wire _temp1289_;
  wire _temp1290_;
  wire _temp1291_;
  wire _temp1292_;
  wire _temp1293_;
  wire _temp1294_;
  wire _temp1295_;
  wire _temp1296_;
  wire _temp1297_;
  wire _temp1298_;
  wire _temp1299_;
  wire _temp1300_;
  wire _temp1301_;
  wire _temp1302_;
  wire _temp1303_;
  wire _temp1304_;
  wire _temp1305_;
  wire _temp1306_;
  wire _temp1307_;
  wire _temp1308_;
  wire _temp1309_;
  wire _temp1310_;
  wire _temp1311_;
  wire _temp1312_;
  wire _temp1313_;
  wire _temp1314_;
  wire _temp1315_;
  wire _temp1316_;
  wire _temp1317_;
  wire _temp1318_;
  wire _temp1319_;
  wire _temp1320_;
  wire _temp1321_;
  wire _temp1322_;
  wire _temp1323_;
  wire _temp1324_;
  wire _temp1325_;
  wire _temp1326_;
  wire _temp1327_;
  wire _temp1328_;
  wire _temp1329_;
  wire _temp1330_;
  wire _temp1331_;
  wire _temp1332_;
  input [31:0] a;
  input [31:0] b;
  output [31:0] q;
  assign _2874_ = b[0] & a[1];
  assign _2885_ = b[1] & a[0];
  assign q[1] = _2885_ ^ _2874_;
  assign q[0] = b[0] & a[0];
  assign _0010_ = b[0] & a[2];
  assign _0021_ = b[1] & a[1];
  assign _0032_ = _0021_ ^ _0010_;
  assign _0043_ = b[2] & a[0];
  assign _temp0_ = _0043_ ^ _0032_;
  assign _0054_ = ~_temp0_;
  assign _0065_ = _2885_ & _2874_;
  assign _0076_ = ~_0065_;
  assign q[2] = _0076_ ^ _0054_;
  assign _0096_ = b[0] & a[3];
  assign _0107_ = b[1] & a[2];
  assign _0118_ = _0107_ ^ _0096_;
  assign _0129_ = b[2] & a[1];
  assign _temp1_ = _0129_ ^ _0118_;
  assign _0140_ = ~_temp1_;
  assign _0151_ = _0021_ & _0010_;
  assign _temp2_ = _0043_ & _0032_;
  assign _temp3_ = _temp2_ | _0151_;
  assign _0162_ = ~_temp3_;
  assign _0173_ = _0162_ ^ _0140_;
  assign _0184_ = b[3] & a[0];
  assign _0194_ = _0184_ ^ _0173_;
  assign _0205_ = _0076_ | _0054_;
  assign _0216_ = ~_0205_;
  assign q[3] = _0216_ ^ _0194_;
  assign _0237_ = b[0] & a[4];
  assign _0248_ = b[1] & a[3];
  assign _0259_ = _0248_ ^ _0237_;
  assign _0270_ = b[2] & a[2];
  assign _temp4_ = _0270_ ^ _0259_;
  assign _0281_ = ~_temp4_;
  assign _0292_ = _0107_ & _0096_;
  assign _temp5_ = _0129_ & _0118_;
  assign _temp6_ = _temp5_ | _0292_;
  assign _0303_ = ~_temp6_;
  assign _0314_ = _0303_ ^ _0281_;
  assign _0324_ = b[3] & a[1];
  assign _0335_ = b[4] & a[0];
  assign _temp7_ = _0335_ ^ _0324_;
  assign _0346_ = ~_temp7_;
  assign _0357_ = _0346_ ^ _0314_;
  assign _temp8_ = _0162_ | _0140_;
  assign _0368_ = ~_temp8_;
  assign _temp9_ = _0184_ & _0173_;
  assign _temp10_ = _temp9_ | _0368_;
  assign _0379_ = ~_temp10_;
  assign _0390_ = _0379_ ^ _0357_;
  assign _0401_ = _0216_ & _0194_;
  assign q[4] = _0401_ ^ _0390_;
  assign _0422_ = b[0] & a[5];
  assign _0433_ = b[1] & a[4];
  assign _0444_ = _0433_ ^ _0422_;
  assign _0454_ = b[2] & a[3];
  assign _temp11_ = _0454_ ^ _0444_;
  assign _0465_ = ~_temp11_;
  assign _0476_ = _0248_ & _0237_;
  assign _temp12_ = _0270_ & _0259_;
  assign _temp13_ = _temp12_ | _0476_;
  assign _0487_ = ~_temp13_;
  assign _0498_ = _0487_ ^ _0465_;
  assign _0509_ = b[3] & a[2];
  assign _0520_ = b[4] & a[1];
  assign _temp14_ = _0520_ ^ _0509_;
  assign _0531_ = ~_temp14_;
  assign _0542_ = b[5] & a[0];
  assign _0553_ = _0542_ ^ _0531_;
  assign _0564_ = _0553_ ^ _0498_;
  assign _0575_ = ~_0346_;
  assign _temp15_ = _0303_ | _0281_;
  assign _0586_ = ~_temp15_;
  assign _temp16_ = _0575_ & _0314_;
  assign _temp17_ = _temp16_ | _0586_;
  assign _0596_ = ~_temp17_;
  assign _0607_ = _0596_ ^ _0564_;
  assign _0618_ = _0335_ & _0324_;
  assign _0629_ = _0618_ ^ _0607_;
  assign _temp18_ = _0379_ | _0357_;
  assign _0640_ = ~_temp18_;
  assign _0651_ = _0640_ ^ _0629_;
  assign _0662_ = _0401_ & _0390_;
  assign q[5] = _0662_ ^ _0651_;
  assign _0683_ = b[0] & a[6];
  assign _0694_ = b[1] & a[5];
  assign _0705_ = _0694_ ^ _0683_;
  assign _0716_ = b[2] & a[4];
  assign _temp19_ = _0716_ ^ _0705_;
  assign _0727_ = ~_temp19_;
  assign _0737_ = _0433_ & _0422_;
  assign _temp20_ = _0454_ & _0444_;
  assign _temp21_ = _temp20_ | _0737_;
  assign _0748_ = ~_temp21_;
  assign _0759_ = _0748_ ^ _0727_;
  assign _0770_ = b[3] & a[3];
  assign _0781_ = b[4] & a[2];
  assign _temp22_ = _0781_ ^ _0770_;
  assign _0792_ = ~_temp22_;
  assign _0803_ = b[5] & a[1];
  assign _0814_ = _0803_ ^ _0792_;
  assign _0825_ = _0814_ ^ _0759_;
  assign _0836_ = ~_0553_;
  assign _temp23_ = _0487_ | _0465_;
  assign _0847_ = ~_temp23_;
  assign _temp24_ = _0836_ & _0498_;
  assign _temp25_ = _temp24_ | _0847_;
  assign _0858_ = ~_temp25_;
  assign _0869_ = _0858_ ^ _0825_;
  assign _0880_ = _0520_ & _0509_;
  assign _0890_ = ~_0531_;
  assign _0901_ = _0542_ & _0890_;
  assign _0912_ = _0901_ | _0880_;
  assign _0923_ = b[6] & a[0];
  assign _0934_ = _0923_ ^ _0912_;
  assign _temp26_ = _0934_ ^ _0869_;
  assign _0945_ = ~_temp26_;
  assign _temp27_ = _0596_ | _0564_;
  assign _0956_ = ~_temp27_;
  assign _temp28_ = _0618_ & _0607_;
  assign _temp29_ = _temp28_ | _0956_;
  assign _0967_ = ~_temp29_;
  assign _0978_ = _0967_ ^ _0945_;
  assign _0989_ = _0640_ & _0629_;
  assign _1000_ = _0989_ ^ _0978_;
  assign _1011_ = _0662_ & _0651_;
  assign q[6] = _1011_ ^ _1000_;
  assign _1032_ = b[0] & a[7];
  assign _1043_ = b[1] & a[6];
  assign _1053_ = _1043_ ^ _1032_;
  assign _1064_ = b[2] & a[5];
  assign _temp30_ = _1064_ ^ _1053_;
  assign _1075_ = ~_temp30_;
  assign _1086_ = _0694_ & _0683_;
  assign _temp31_ = _0716_ & _0705_;
  assign _temp32_ = _temp31_ | _1086_;
  assign _1097_ = ~_temp32_;
  assign _1108_ = _1097_ ^ _1075_;
  assign _1119_ = b[3] & a[4];
  assign _1130_ = b[4] & a[3];
  assign _1141_ = _1130_ ^ _1119_;
  assign _1152_ = b[5] & a[2];
  assign _1163_ = _1152_ ^ _1141_;
  assign _temp33_ = _1163_ ^ _1108_;
  assign _1174_ = ~_temp33_;
  assign _1185_ = ~_0814_;
  assign _temp34_ = _0748_ | _0727_;
  assign _1196_ = ~_temp34_;
  assign _temp35_ = _1185_ & _0759_;
  assign _temp36_ = _temp35_ | _1196_;
  assign _1207_ = ~_temp36_;
  assign _1218_ = _1207_ ^ _1174_;
  assign _1228_ = _0781_ & _0770_;
  assign _1239_ = ~_0792_;
  assign _1250_ = _0803_ & _1239_;
  assign _temp37_ = _1250_ | _1228_;
  assign _1261_ = ~_temp37_;
  assign _1272_ = b[6] & a[1];
  assign _1283_ = b[7] & a[0];
  assign _temp38_ = _1283_ ^ _1272_;
  assign _1294_ = ~_temp38_;
  assign _1305_ = _1294_ ^ _1261_;
  assign _temp39_ = _1305_ ^ _1218_;
  assign _1316_ = ~_temp39_;
  assign _temp40_ = _0858_ | _0825_;
  assign _1327_ = ~_temp40_;
  assign _temp41_ = _0934_ & _0869_;
  assign _temp42_ = _temp41_ | _1327_;
  assign _1338_ = ~_temp42_;
  assign _1349_ = _1338_ ^ _1316_;
  assign _1360_ = _0923_ & _0912_;
  assign _1371_ = _1360_ ^ _1349_;
  assign _temp43_ = _0967_ | _0945_;
  assign _1382_ = ~_temp43_;
  assign _1393_ = _1382_ ^ _1371_;
  assign _1404_ = _0989_ & _0978_;
  assign _1414_ = _1404_ ^ _1393_;
  assign _1425_ = _1011_ & _1000_;
  assign q[7] = _1425_ ^ _1414_;
  assign _1446_ = a[8] & b[0];
  assign _1457_ = b[1] & a[7];
  assign _1468_ = _1457_ ^ _1446_;
  assign _1479_ = b[2] & a[6];
  assign _temp44_ = _1479_ ^ _1468_;
  assign _1490_ = ~_temp44_;
  assign _1501_ = _1043_ & _1032_;
  assign _temp45_ = _1064_ & _1053_;
  assign _temp46_ = _temp45_ | _1501_;
  assign _1512_ = ~_temp46_;
  assign _1523_ = _1512_ ^ _1490_;
  assign _1534_ = b[3] & a[5];
  assign _1545_ = b[4] & a[4];
  assign _1556_ = _1545_ ^ _1534_;
  assign _1567_ = b[5] & a[3];
  assign _1578_ = _1567_ ^ _1556_;
  assign _temp47_ = _1578_ ^ _1523_;
  assign _1589_ = ~_temp47_;
  assign _temp48_ = _1097_ | _1075_;
  assign _1600_ = ~_temp48_;
  assign _temp49_ = _1163_ & _1108_;
  assign _temp50_ = _temp49_ | _1600_;
  assign _1611_ = ~_temp50_;
  assign _1621_ = _1611_ ^ _1589_;
  assign _1632_ = _1130_ & _1119_;
  assign _1643_ = _1152_ & _1141_;
  assign _temp51_ = _1643_ | _1632_;
  assign _1654_ = ~_temp51_;
  assign _1665_ = b[6] & a[2];
  assign _1676_ = b[7] & a[1];
  assign _1687_ = _1676_ ^ _1665_;
  assign _1698_ = b[8] & a[0];
  assign _temp52_ = _1698_ ^ _1687_;
  assign _1709_ = ~_temp52_;
  assign _1720_ = _1709_ ^ _1654_;
  assign _1731_ = _1283_ & _1272_;
  assign _1742_ = _1731_ ^ _1720_;
  assign _temp53_ = _1742_ ^ _1621_;
  assign _1753_ = ~_temp53_;
  assign _temp54_ = _1207_ | _1174_;
  assign _1764_ = ~_temp54_;
  assign _temp55_ = _1305_ & _1218_;
  assign _temp56_ = _temp55_ | _1764_;
  assign _1775_ = ~_temp56_;
  assign _1786_ = _1775_ ^ _1753_;
  assign _temp57_ = _1294_ | _1261_;
  assign _1797_ = ~_temp57_;
  assign _temp58_ = _1797_ ^ _1786_;
  assign _1808_ = ~_temp58_;
  assign _temp59_ = _1338_ | _1316_;
  assign _1818_ = ~_temp59_;
  assign _temp60_ = _1360_ & _1349_;
  assign _temp61_ = _temp60_ | _1818_;
  assign _1829_ = ~_temp61_;
  assign _1840_ = _1829_ ^ _1808_;
  assign _1851_ = _1382_ & _1371_;
  assign _1862_ = _1851_ ^ _1840_;
  assign _1873_ = _1404_ & _1393_;
  assign _1884_ = _1873_ ^ _1862_;
  assign _1895_ = _1425_ & _1414_;
  assign q[8] = _1895_ ^ _1884_;
  assign _1916_ = a[9] & b[0];
  assign _1927_ = b[1] & a[8];
  assign _1938_ = _1927_ ^ _1916_;
  assign _1949_ = b[2] & a[7];
  assign _temp62_ = _1949_ ^ _1938_;
  assign _1960_ = ~_temp62_;
  assign _1971_ = _1457_ & _1446_;
  assign _temp63_ = _1479_ & _1468_;
  assign _temp64_ = _temp63_ | _1971_;
  assign _1982_ = ~_temp64_;
  assign _1993_ = _1982_ ^ _1960_;
  assign _2004_ = b[3] & a[6];
  assign _2015_ = b[4] & a[5];
  assign _2025_ = _2015_ ^ _2004_;
  assign _2046_ = b[5] & a[4];
  assign _2047_ = _2046_ ^ _2025_;
  assign _temp65_ = _2047_ ^ _1993_;
  assign _2058_ = ~_temp65_;
  assign _temp66_ = _1512_ | _1490_;
  assign _2069_ = ~_temp66_;
  assign _temp67_ = _1578_ & _1523_;
  assign _temp68_ = _temp67_ | _2069_;
  assign _2080_ = ~_temp68_;
  assign _2091_ = _2080_ ^ _2058_;
  assign _2102_ = _1545_ & _1534_;
  assign _2113_ = _1567_ & _1556_;
  assign _temp69_ = _2113_ | _2102_;
  assign _2124_ = ~_temp69_;
  assign _2135_ = b[6] & a[3];
  assign _2146_ = b[7] & a[2];
  assign _2157_ = _2146_ ^ _2135_;
  assign _2168_ = b[8] & a[1];
  assign _temp70_ = _2168_ ^ _2157_;
  assign _2179_ = ~_temp70_;
  assign _2190_ = _2179_ ^ _2124_;
  assign _2201_ = _1676_ & _1665_;
  assign _2212_ = _1698_ & _1687_;
  assign _2217_ = _2212_ | _2201_;
  assign _2218_ = _2217_ ^ _2190_;
  assign _temp71_ = _2218_ ^ _2091_;
  assign _2219_ = ~_temp71_;
  assign _temp72_ = _1611_ | _1589_;
  assign _2220_ = ~_temp72_;
  assign _temp73_ = _1742_ & _1621_;
  assign _temp74_ = _temp73_ | _2220_;
  assign _2221_ = ~_temp74_;
  assign _2222_ = _2221_ ^ _2219_;
  assign _temp75_ = _1709_ | _1654_;
  assign _2223_ = ~_temp75_;
  assign _2224_ = _1731_ & _1720_;
  assign _2225_ = _2224_ | _2223_;
  assign _2226_ = b[9] & a[0];
  assign _2227_ = _2226_ ^ _2225_;
  assign _temp76_ = _2227_ ^ _2222_;
  assign _2228_ = ~_temp76_;
  assign _temp77_ = _1775_ | _1753_;
  assign _2229_ = ~_temp77_;
  assign _temp78_ = _1797_ & _1786_;
  assign _temp79_ = _temp78_ | _2229_;
  assign _2230_ = ~_temp79_;
  assign _2231_ = _2230_ ^ _2228_;
  assign _temp80_ = _1829_ | _1808_;
  assign _2232_ = ~_temp80_;
  assign _2233_ = _2232_ ^ _2231_;
  assign _2234_ = _1851_ & _1840_;
  assign _2235_ = _2234_ ^ _2233_;
  assign _2236_ = _1873_ & _1862_;
  assign _2237_ = _2236_ ^ _2235_;
  assign _2238_ = _1895_ & _1884_;
  assign q[9] = _2238_ ^ _2237_;
  assign _2239_ = a[10] & b[0];
  assign _2240_ = b[1] & a[9];
  assign _2241_ = _2240_ ^ _2239_;
  assign _2242_ = b[2] & a[8];
  assign _temp81_ = _2242_ ^ _2241_;
  assign _2243_ = ~_temp81_;
  assign _2244_ = _1927_ & _1916_;
  assign _temp82_ = _1949_ & _1938_;
  assign _temp83_ = _temp82_ | _2244_;
  assign _2245_ = ~_temp83_;
  assign _2246_ = _2245_ ^ _2243_;
  assign _2247_ = b[3] & a[7];
  assign _2248_ = b[4] & a[6];
  assign _2249_ = _2248_ ^ _2247_;
  assign _2250_ = b[5] & a[5];
  assign _2251_ = _2250_ ^ _2249_;
  assign _temp84_ = _2251_ ^ _2246_;
  assign _2252_ = ~_temp84_;
  assign _temp85_ = _1982_ | _1960_;
  assign _2253_ = ~_temp85_;
  assign _temp86_ = _2047_ & _1993_;
  assign _temp87_ = _temp86_ | _2253_;
  assign _2254_ = ~_temp87_;
  assign _2255_ = _2254_ ^ _2252_;
  assign _2256_ = _2015_ & _2004_;
  assign _2257_ = _2046_ & _2025_;
  assign _temp88_ = _2257_ | _2256_;
  assign _2258_ = ~_temp88_;
  assign _2259_ = b[6] & a[4];
  assign _2260_ = b[7] & a[3];
  assign _2261_ = _2260_ ^ _2259_;
  assign _2262_ = b[8] & a[2];
  assign _temp89_ = _2262_ ^ _2261_;
  assign _2263_ = ~_temp89_;
  assign _2264_ = _2263_ ^ _2258_;
  assign _2265_ = _2146_ & _2135_;
  assign _2266_ = _2168_ & _2157_;
  assign _2267_ = _2266_ | _2265_;
  assign _2268_ = _2267_ ^ _2264_;
  assign _temp90_ = _2268_ ^ _2255_;
  assign _2269_ = ~_temp90_;
  assign _temp91_ = _2080_ | _2058_;
  assign _2270_ = ~_temp91_;
  assign _temp92_ = _2218_ & _2091_;
  assign _temp93_ = _temp92_ | _2270_;
  assign _2271_ = ~_temp93_;
  assign _2272_ = _2271_ ^ _2269_;
  assign _temp94_ = _2179_ | _2124_;
  assign _2273_ = ~_temp94_;
  assign _2274_ = _2217_ & _2190_;
  assign _temp95_ = _2274_ | _2273_;
  assign _2275_ = ~_temp95_;
  assign _2276_ = b[9] & a[1];
  assign _2277_ = b[10] & a[0];
  assign _temp96_ = _2277_ ^ _2276_;
  assign _2278_ = ~_temp96_;
  assign _2279_ = _2278_ ^ _2275_;
  assign _temp97_ = _2279_ ^ _2272_;
  assign _2280_ = ~_temp97_;
  assign _temp98_ = _2221_ | _2219_;
  assign _2281_ = ~_temp98_;
  assign _temp99_ = _2227_ & _2222_;
  assign _temp100_ = _temp99_ | _2281_;
  assign _2282_ = ~_temp100_;
  assign _2283_ = _2282_ ^ _2280_;
  assign _2284_ = _2226_ & _2225_;
  assign _2285_ = _2284_ ^ _2283_;
  assign _temp101_ = _2230_ | _2228_;
  assign _2286_ = ~_temp101_;
  assign _2287_ = _2286_ ^ _2285_;
  assign _2288_ = _2232_ & _2231_;
  assign _2289_ = _2288_ ^ _2287_;
  assign _2290_ = _2234_ & _2233_;
  assign _2291_ = _2290_ ^ _2289_;
  assign _2292_ = _2236_ & _2235_;
  assign _2293_ = _2292_ ^ _2291_;
  assign _2294_ = _2238_ & _2237_;
  assign q[10] = _2294_ ^ _2293_;
  assign _2295_ = a[11] & b[0];
  assign _2296_ = b[1] & a[10];
  assign _2297_ = _2296_ ^ _2295_;
  assign _2298_ = b[2] & a[9];
  assign _temp102_ = _2298_ ^ _2297_;
  assign _2299_ = ~_temp102_;
  assign _2300_ = _2240_ & _2239_;
  assign _temp103_ = _2242_ & _2241_;
  assign _temp104_ = _temp103_ | _2300_;
  assign _2301_ = ~_temp104_;
  assign _2302_ = _2301_ ^ _2299_;
  assign _2303_ = b[3] & a[8];
  assign _2304_ = b[4] & a[7];
  assign _2305_ = _2304_ ^ _2303_;
  assign _2306_ = b[5] & a[6];
  assign _2307_ = _2306_ ^ _2305_;
  assign _temp105_ = _2307_ ^ _2302_;
  assign _2308_ = ~_temp105_;
  assign _temp106_ = _2245_ | _2243_;
  assign _2309_ = ~_temp106_;
  assign _temp107_ = _2251_ & _2246_;
  assign _temp108_ = _temp107_ | _2309_;
  assign _2310_ = ~_temp108_;
  assign _2311_ = _2310_ ^ _2308_;
  assign _2312_ = _2248_ & _2247_;
  assign _2313_ = _2250_ & _2249_;
  assign _temp109_ = _2313_ | _2312_;
  assign _2314_ = ~_temp109_;
  assign _2315_ = b[6] & a[5];
  assign _2316_ = b[7] & a[4];
  assign _2317_ = _2316_ ^ _2315_;
  assign _2318_ = b[8] & a[3];
  assign _temp110_ = _2318_ ^ _2317_;
  assign _2319_ = ~_temp110_;
  assign _2320_ = _2319_ ^ _2314_;
  assign _2321_ = _2260_ & _2259_;
  assign _2322_ = _2262_ & _2261_;
  assign _2323_ = _2322_ | _2321_;
  assign _2324_ = _2323_ ^ _2320_;
  assign _temp111_ = _2324_ ^ _2311_;
  assign _2325_ = ~_temp111_;
  assign _temp112_ = _2254_ | _2252_;
  assign _2326_ = ~_temp112_;
  assign _temp113_ = _2268_ & _2255_;
  assign _temp114_ = _temp113_ | _2326_;
  assign _2327_ = ~_temp114_;
  assign _2328_ = _2327_ ^ _2325_;
  assign _temp115_ = _2263_ | _2258_;
  assign _2329_ = ~_temp115_;
  assign _2330_ = _2267_ & _2264_;
  assign _temp116_ = _2330_ | _2329_;
  assign _2331_ = ~_temp116_;
  assign _2332_ = b[9] & a[2];
  assign _2333_ = b[10] & a[1];
  assign _2334_ = _2333_ ^ _2332_;
  assign _2335_ = b[11] & a[0];
  assign _temp117_ = _2335_ ^ _2334_;
  assign _2336_ = ~_temp117_;
  assign _2337_ = _2277_ & _2276_;
  assign _2338_ = _2337_ ^ _2336_;
  assign _2339_ = _2338_ ^ _2331_;
  assign _temp118_ = _2339_ ^ _2328_;
  assign _2340_ = ~_temp118_;
  assign _temp119_ = _2271_ | _2269_;
  assign _2341_ = ~_temp119_;
  assign _temp120_ = _2279_ & _2272_;
  assign _temp121_ = _temp120_ | _2341_;
  assign _2342_ = ~_temp121_;
  assign _2343_ = _2342_ ^ _2340_;
  assign _temp122_ = _2278_ | _2275_;
  assign _2344_ = ~_temp122_;
  assign _temp123_ = _2344_ ^ _2343_;
  assign _2345_ = ~_temp123_;
  assign _temp124_ = _2282_ | _2280_;
  assign _2346_ = ~_temp124_;
  assign _temp125_ = _2284_ & _2283_;
  assign _temp126_ = _temp125_ | _2346_;
  assign _2347_ = ~_temp126_;
  assign _2348_ = _2347_ ^ _2345_;
  assign _2349_ = _2286_ & _2285_;
  assign _2350_ = _2349_ ^ _2348_;
  assign _2351_ = _2288_ & _2287_;
  assign _2352_ = _2351_ ^ _2350_;
  assign _2353_ = _2290_ & _2289_;
  assign _temp127_ = _2353_ ^ _2352_;
  assign _2354_ = ~_temp127_;
  assign _2355_ = _2292_ & _2291_;
  assign _temp128_ = _2294_ & _2293_;
  assign _temp129_ = _temp128_ | _2355_;
  assign _2356_ = ~_temp129_;
  assign q[11] = _2356_ ^ _2354_;
  assign _2357_ = a[12] & b[0];
  assign _2358_ = b[1] & a[11];
  assign _2359_ = _2358_ ^ _2357_;
  assign _2360_ = b[2] & a[10];
  assign _temp130_ = _2360_ ^ _2359_;
  assign _2361_ = ~_temp130_;
  assign _2362_ = _2296_ & _2295_;
  assign _temp131_ = _2298_ & _2297_;
  assign _temp132_ = _temp131_ | _2362_;
  assign _2363_ = ~_temp132_;
  assign _2364_ = _2363_ ^ _2361_;
  assign _2365_ = b[3] & a[9];
  assign _2366_ = b[4] & a[8];
  assign _2367_ = _2366_ ^ _2365_;
  assign _2368_ = b[5] & a[7];
  assign _2369_ = _2368_ ^ _2367_;
  assign _temp133_ = _2369_ ^ _2364_;
  assign _2370_ = ~_temp133_;
  assign _temp134_ = _2301_ | _2299_;
  assign _2371_ = ~_temp134_;
  assign _temp135_ = _2307_ & _2302_;
  assign _temp136_ = _temp135_ | _2371_;
  assign _2372_ = ~_temp136_;
  assign _2373_ = _2372_ ^ _2370_;
  assign _2374_ = _2304_ & _2303_;
  assign _2375_ = _2306_ & _2305_;
  assign _temp137_ = _2375_ | _2374_;
  assign _2376_ = ~_temp137_;
  assign _2377_ = b[6] & a[6];
  assign _2378_ = b[7] & a[5];
  assign _2379_ = _2378_ ^ _2377_;
  assign _2380_ = b[8] & a[4];
  assign _temp138_ = _2380_ ^ _2379_;
  assign _2381_ = ~_temp138_;
  assign _temp139_ = _2381_ ^ _2376_;
  assign _2382_ = ~_temp139_;
  assign _2383_ = _2316_ & _2315_;
  assign _2384_ = _2318_ & _2317_;
  assign _temp140_ = _2384_ | _2383_;
  assign _2385_ = ~_temp140_;
  assign _2386_ = _2385_ ^ _2382_;
  assign _temp141_ = _2386_ ^ _2373_;
  assign _2387_ = ~_temp141_;
  assign _temp142_ = _2310_ | _2308_;
  assign _2388_ = ~_temp142_;
  assign _temp143_ = _2324_ & _2311_;
  assign _temp144_ = _temp143_ | _2388_;
  assign _2389_ = ~_temp144_;
  assign _2390_ = _2389_ ^ _2387_;
  assign _temp145_ = _2319_ | _2314_;
  assign _2391_ = ~_temp145_;
  assign _2392_ = _2323_ & _2320_;
  assign _temp146_ = _2392_ | _2391_;
  assign _2393_ = ~_temp146_;
  assign _2394_ = b[9] & a[3];
  assign _2395_ = b[10] & a[2];
  assign _2396_ = _2395_ ^ _2394_;
  assign _2397_ = b[11] & a[1];
  assign _temp147_ = _2397_ ^ _2396_;
  assign _2398_ = ~_temp147_;
  assign _2399_ = _2333_ & _2332_;
  assign _temp148_ = _2335_ & _2334_;
  assign _temp149_ = _temp148_ | _2399_;
  assign _2400_ = ~_temp149_;
  assign _2401_ = _2400_ ^ _2398_;
  assign _2402_ = b[12] & a[0];
  assign _temp150_ = _2402_ ^ _2401_;
  assign _2403_ = ~_temp150_;
  assign _2404_ = _2403_ ^ _2393_;
  assign _2405_ = ~_2337_;
  assign _temp151_ = _2405_ | _2336_;
  assign _2406_ = ~_temp151_;
  assign _2407_ = _2406_ ^ _2404_;
  assign _temp152_ = _2407_ ^ _2390_;
  assign _2408_ = ~_temp152_;
  assign _temp153_ = _2327_ | _2325_;
  assign _2409_ = ~_temp153_;
  assign _temp154_ = _2339_ & _2328_;
  assign _temp155_ = _temp154_ | _2409_;
  assign _2410_ = ~_temp155_;
  assign _2411_ = _2410_ ^ _2408_;
  assign _temp156_ = _2338_ | _2331_;
  assign _2412_ = ~_temp156_;
  assign _temp157_ = _2412_ ^ _2411_;
  assign _2413_ = ~_temp157_;
  assign _temp158_ = _2342_ | _2340_;
  assign _2414_ = ~_temp158_;
  assign _temp159_ = _2344_ & _2343_;
  assign _temp160_ = _temp159_ | _2414_;
  assign _2415_ = ~_temp160_;
  assign _2416_ = _2415_ ^ _2413_;
  assign _temp161_ = _2347_ | _2345_;
  assign _2417_ = ~_temp161_;
  assign _2418_ = _2417_ ^ _2416_;
  assign _2419_ = _2349_ & _2348_;
  assign _2420_ = _2419_ ^ _2418_;
  assign _2421_ = _2351_ & _2350_;
  assign _2422_ = _2421_ ^ _2420_;
  assign _temp162_ = _2294_ & _2293_;
  assign _2423_ = ~_temp162_;
  assign _2424_ = _2353_ ^ _2352_;
  assign _2425_ = _2353_ & _2352_;
  assign _temp163_ = _2355_ & _2424_;
  assign _temp164_ = _temp163_ | _2425_;
  assign _2426_ = ~_temp164_;
  assign _temp165_ = _2423_ | _2354_;
  assign _temp166_ = _temp165_ & _2426_;
  assign _2427_ = ~_temp166_;
  assign q[12] = _2427_ ^ _2422_;
  assign _2428_ = a[13] & b[0];
  assign _2429_ = b[1] & a[12];
  assign _2430_ = _2429_ ^ _2428_;
  assign _2431_ = b[2] & a[11];
  assign _temp167_ = _2431_ ^ _2430_;
  assign _2432_ = ~_temp167_;
  assign _2433_ = _2358_ & _2357_;
  assign _temp168_ = _2360_ & _2359_;
  assign _temp169_ = _temp168_ | _2433_;
  assign _2434_ = ~_temp169_;
  assign _2435_ = _2434_ ^ _2432_;
  assign _2436_ = b[3] & a[10];
  assign _2437_ = b[4] & a[9];
  assign _2438_ = _2437_ ^ _2436_;
  assign _2439_ = b[5] & a[8];
  assign _2440_ = _2439_ ^ _2438_;
  assign _temp170_ = _2440_ ^ _2435_;
  assign _2441_ = ~_temp170_;
  assign _temp171_ = _2363_ | _2361_;
  assign _2442_ = ~_temp171_;
  assign _temp172_ = _2369_ & _2364_;
  assign _temp173_ = _temp172_ | _2442_;
  assign _2443_ = ~_temp173_;
  assign _2444_ = _2443_ ^ _2441_;
  assign _2445_ = _2366_ & _2365_;
  assign _2446_ = _2368_ & _2367_;
  assign _temp174_ = _2446_ | _2445_;
  assign _2447_ = ~_temp174_;
  assign _2448_ = b[6] & a[7];
  assign _2449_ = b[7] & a[6];
  assign _2450_ = _2449_ ^ _2448_;
  assign _2451_ = b[8] & a[5];
  assign _temp175_ = _2451_ ^ _2450_;
  assign _2452_ = ~_temp175_;
  assign _temp176_ = _2452_ ^ _2447_;
  assign _2453_ = ~_temp176_;
  assign _2454_ = _2378_ & _2377_;
  assign _2455_ = _2380_ & _2379_;
  assign _temp177_ = _2455_ | _2454_;
  assign _2456_ = ~_temp177_;
  assign _2457_ = _2456_ ^ _2453_;
  assign _temp178_ = _2457_ ^ _2444_;
  assign _2458_ = ~_temp178_;
  assign _temp179_ = _2372_ | _2370_;
  assign _2459_ = ~_temp179_;
  assign _temp180_ = _2386_ & _2373_;
  assign _temp181_ = _temp180_ | _2459_;
  assign _2460_ = ~_temp181_;
  assign _2461_ = _2460_ ^ _2458_;
  assign _2462_ = _2381_ ^ _2376_;
  assign _2463_ = _2384_ | _2383_;
  assign _temp182_ = _2381_ | _2376_;
  assign _2464_ = ~_temp182_;
  assign _temp183_ = _2463_ & _2462_;
  assign _temp184_ = _temp183_ | _2464_;
  assign _2465_ = ~_temp184_;
  assign _2466_ = b[9] & a[4];
  assign _2467_ = b[10] & a[3];
  assign _2468_ = _2467_ ^ _2466_;
  assign _2469_ = b[11] & a[2];
  assign _temp185_ = _2469_ ^ _2468_;
  assign _2470_ = ~_temp185_;
  assign _2471_ = _2395_ & _2394_;
  assign _temp186_ = _2397_ & _2396_;
  assign _temp187_ = _temp186_ | _2471_;
  assign _2472_ = ~_temp187_;
  assign _2473_ = _2472_ ^ _2470_;
  assign _2474_ = b[12] & a[1];
  assign _2475_ = b[13] & a[0];
  assign _temp188_ = _2475_ ^ _2474_;
  assign _2476_ = ~_temp188_;
  assign _2477_ = _2476_ ^ _2473_;
  assign _2478_ = _2477_ ^ _2465_;
  assign _temp189_ = _2400_ | _2398_;
  assign _2479_ = ~_temp189_;
  assign _2480_ = _2402_ & _2401_;
  assign _2481_ = _2480_ | _2479_;
  assign _2482_ = _2481_ ^ _2478_;
  assign _temp190_ = _2482_ ^ _2461_;
  assign _2483_ = ~_temp190_;
  assign _temp191_ = _2389_ | _2387_;
  assign _2484_ = ~_temp191_;
  assign _temp192_ = _2407_ & _2390_;
  assign _temp193_ = _temp192_ | _2484_;
  assign _2485_ = ~_temp193_;
  assign _2486_ = _2485_ ^ _2483_;
  assign _temp194_ = _2403_ | _2393_;
  assign _2487_ = ~_temp194_;
  assign _2488_ = _2406_ & _2404_;
  assign _temp195_ = _2488_ | _2487_;
  assign _2489_ = ~_temp195_;
  assign _2490_ = _2489_ ^ _2486_;
  assign _temp196_ = _2410_ | _2408_;
  assign _2491_ = ~_temp196_;
  assign _temp197_ = _2412_ & _2411_;
  assign _temp198_ = _temp197_ | _2491_;
  assign _2492_ = ~_temp198_;
  assign _2493_ = _2492_ ^ _2490_;
  assign _temp199_ = _2415_ | _2413_;
  assign _2494_ = ~_temp199_;
  assign _2495_ = _2494_ ^ _2493_;
  assign _2496_ = _2417_ & _2416_;
  assign _2497_ = _2496_ ^ _2495_;
  assign _2498_ = _2419_ & _2418_;
  assign _2499_ = _2498_ ^ _2497_;
  assign _2500_ = _2421_ & _2420_;
  assign _temp200_ = _2427_ & _2422_;
  assign _temp201_ = _temp200_ | _2500_;
  assign _2501_ = ~_temp201_;
  assign _temp202_ = _2501_ ^ _2499_;
  assign q[13] = ~_temp202_;
  assign _2502_ = a[14] & b[0];
  assign _2503_ = b[1] & a[13];
  assign _2504_ = _2503_ ^ _2502_;
  assign _2505_ = b[2] & a[12];
  assign _temp203_ = _2505_ ^ _2504_;
  assign _2506_ = ~_temp203_;
  assign _2507_ = _2429_ & _2428_;
  assign _temp204_ = _2431_ & _2430_;
  assign _temp205_ = _temp204_ | _2507_;
  assign _2508_ = ~_temp205_;
  assign _2509_ = _2508_ ^ _2506_;
  assign _2510_ = b[3] & a[11];
  assign _2511_ = b[4] & a[10];
  assign _2512_ = _2511_ ^ _2510_;
  assign _2513_ = b[5] & a[9];
  assign _2514_ = _2513_ ^ _2512_;
  assign _temp206_ = _2514_ ^ _2509_;
  assign _2515_ = ~_temp206_;
  assign _temp207_ = _2434_ | _2432_;
  assign _2516_ = ~_temp207_;
  assign _temp208_ = _2440_ & _2435_;
  assign _temp209_ = _temp208_ | _2516_;
  assign _2517_ = ~_temp209_;
  assign _2518_ = _2517_ ^ _2515_;
  assign _2519_ = _2437_ & _2436_;
  assign _2520_ = _2439_ & _2438_;
  assign _temp210_ = _2520_ | _2519_;
  assign _2521_ = ~_temp210_;
  assign _2522_ = b[6] & a[8];
  assign _2523_ = b[7] & a[7];
  assign _2524_ = _2523_ ^ _2522_;
  assign _2525_ = b[8] & a[6];
  assign _temp211_ = _2525_ ^ _2524_;
  assign _2526_ = ~_temp211_;
  assign _2527_ = _2526_ ^ _2521_;
  assign _2528_ = _2449_ & _2448_;
  assign _2529_ = _2451_ & _2450_;
  assign _2530_ = _2529_ | _2528_;
  assign _2531_ = _2530_ ^ _2527_;
  assign _temp212_ = _2531_ ^ _2518_;
  assign _2532_ = ~_temp212_;
  assign _temp213_ = _2443_ | _2441_;
  assign _2533_ = ~_temp213_;
  assign _temp214_ = _2457_ & _2444_;
  assign _temp215_ = _temp214_ | _2533_;
  assign _2534_ = ~_temp215_;
  assign _2535_ = _2534_ ^ _2532_;
  assign _2536_ = _2452_ ^ _2447_;
  assign _2537_ = _2455_ | _2454_;
  assign _temp216_ = _2452_ | _2447_;
  assign _2538_ = ~_temp216_;
  assign _temp217_ = _2537_ & _2536_;
  assign _temp218_ = _temp217_ | _2538_;
  assign _2539_ = ~_temp218_;
  assign _2540_ = b[9] & a[5];
  assign _2541_ = b[10] & a[4];
  assign _2542_ = _2541_ ^ _2540_;
  assign _2543_ = b[11] & a[3];
  assign _temp219_ = _2543_ ^ _2542_;
  assign _2544_ = ~_temp219_;
  assign _2545_ = _2467_ & _2466_;
  assign _temp220_ = _2469_ & _2468_;
  assign _temp221_ = _temp220_ | _2545_;
  assign _2546_ = ~_temp221_;
  assign _2547_ = _2546_ ^ _2544_;
  assign _2548_ = b[12] & a[2];
  assign _2549_ = b[13] & a[1];
  assign _temp222_ = _2549_ ^ _2548_;
  assign _2550_ = ~_temp222_;
  assign _2551_ = b[14] & a[0];
  assign _2552_ = _2551_ ^ _2550_;
  assign _2553_ = _2552_ ^ _2547_;
  assign _2554_ = _2553_ ^ _2539_;
  assign _temp223_ = _2472_ | _2470_;
  assign _2555_ = ~_temp223_;
  assign _2556_ = ~_2476_;
  assign _2557_ = _2556_ & _2473_;
  assign _2558_ = _2557_ | _2555_;
  assign _2559_ = _2558_ ^ _2554_;
  assign _temp224_ = _2559_ ^ _2535_;
  assign _2560_ = ~_temp224_;
  assign _temp225_ = _2460_ | _2458_;
  assign _2561_ = ~_temp225_;
  assign _temp226_ = _2482_ & _2461_;
  assign _temp227_ = _temp226_ | _2561_;
  assign _2562_ = ~_temp227_;
  assign _2563_ = _2562_ ^ _2560_;
  assign _temp228_ = _2477_ | _2465_;
  assign _2564_ = ~_temp228_;
  assign _2565_ = _2481_ & _2478_;
  assign _2566_ = _2565_ | _2564_;
  assign _2567_ = _2475_ & _2474_;
  assign _2568_ = _2567_ ^ _2566_;
  assign _temp229_ = _2568_ ^ _2563_;
  assign _2569_ = ~_temp229_;
  assign _2570_ = ~_2489_;
  assign _temp230_ = _2485_ | _2483_;
  assign _2571_ = ~_temp230_;
  assign _temp231_ = _2570_ & _2486_;
  assign _temp232_ = _temp231_ | _2571_;
  assign _2572_ = ~_temp232_;
  assign _2573_ = _2572_ ^ _2569_;
  assign _temp233_ = _2492_ | _2490_;
  assign _2574_ = ~_temp233_;
  assign _2575_ = _2574_ ^ _2573_;
  assign _2576_ = _2494_ & _2493_;
  assign _2577_ = _2576_ ^ _2575_;
  assign _2578_ = _2496_ & _2495_;
  assign _2579_ = _2578_ ^ _2577_;
  assign _2580_ = _2498_ & _2497_;
  assign _2581_ = _2500_ & _2499_;
  assign _temp234_ = _2581_ | _2580_;
  assign _2582_ = ~_temp234_;
  assign _2583_ = ~_2582_;
  assign _2584_ = _2499_ & _2422_;
  assign _2585_ = _2584_ & _2427_;
  assign _2586_ = _2585_ | _2583_;
  assign q[14] = _2586_ ^ _2579_;
  assign _2587_ = a[15] & b[0];
  assign _2588_ = b[1] & a[14];
  assign _2589_ = _2588_ ^ _2587_;
  assign _2590_ = b[2] & a[13];
  assign _temp235_ = _2590_ ^ _2589_;
  assign _2591_ = ~_temp235_;
  assign _2592_ = _2503_ & _2502_;
  assign _temp236_ = _2505_ & _2504_;
  assign _temp237_ = _temp236_ | _2592_;
  assign _2593_ = ~_temp237_;
  assign _2594_ = _2593_ ^ _2591_;
  assign _2595_ = b[3] & a[12];
  assign _2596_ = b[4] & a[11];
  assign _2597_ = _2596_ ^ _2595_;
  assign _2598_ = b[5] & a[10];
  assign _2599_ = _2598_ ^ _2597_;
  assign _temp238_ = _2599_ ^ _2594_;
  assign _2600_ = ~_temp238_;
  assign _temp239_ = _2508_ | _2506_;
  assign _2601_ = ~_temp239_;
  assign _temp240_ = _2514_ & _2509_;
  assign _temp241_ = _temp240_ | _2601_;
  assign _2602_ = ~_temp241_;
  assign _2603_ = _2602_ ^ _2600_;
  assign _2604_ = _2511_ & _2510_;
  assign _2605_ = _2513_ & _2512_;
  assign _temp242_ = _2605_ | _2604_;
  assign _2606_ = ~_temp242_;
  assign _2607_ = b[6] & a[9];
  assign _2608_ = b[7] & a[8];
  assign _2609_ = _2608_ ^ _2607_;
  assign _2610_ = b[8] & a[7];
  assign _temp243_ = _2610_ ^ _2609_;
  assign _2611_ = ~_temp243_;
  assign _2612_ = _2611_ ^ _2606_;
  assign _2613_ = _2523_ & _2522_;
  assign _2614_ = _2525_ & _2524_;
  assign _2615_ = _2614_ | _2613_;
  assign _2616_ = _2615_ ^ _2612_;
  assign _temp244_ = _2616_ ^ _2603_;
  assign _2617_ = ~_temp244_;
  assign _temp245_ = _2517_ | _2515_;
  assign _2618_ = ~_temp245_;
  assign _temp246_ = _2531_ & _2518_;
  assign _temp247_ = _temp246_ | _2618_;
  assign _2619_ = ~_temp247_;
  assign _2620_ = _2619_ ^ _2617_;
  assign _temp248_ = _2526_ | _2521_;
  assign _2621_ = ~_temp248_;
  assign _temp249_ = _2530_ & _2527_;
  assign _temp250_ = _temp249_ | _2621_;
  assign _2622_ = ~_temp250_;
  assign _2623_ = b[9] & a[6];
  assign _2624_ = b[10] & a[5];
  assign _2625_ = _2624_ ^ _2623_;
  assign _2626_ = b[11] & a[4];
  assign _temp251_ = _2626_ ^ _2625_;
  assign _2627_ = ~_temp251_;
  assign _2628_ = _2541_ & _2540_;
  assign _temp252_ = _2543_ & _2542_;
  assign _temp253_ = _temp252_ | _2628_;
  assign _2629_ = ~_temp253_;
  assign _2630_ = _2629_ ^ _2627_;
  assign _2631_ = b[12] & a[3];
  assign _2632_ = b[13] & a[2];
  assign _temp254_ = _2632_ ^ _2631_;
  assign _2633_ = ~_temp254_;
  assign _2634_ = b[14] & a[1];
  assign _2635_ = _2634_ ^ _2633_;
  assign _2636_ = _2635_ ^ _2630_;
  assign _2637_ = _2636_ ^ _2622_;
  assign _temp255_ = _2546_ | _2544_;
  assign _2638_ = ~_temp255_;
  assign _2639_ = ~_2552_;
  assign _2640_ = _2639_ & _2547_;
  assign _temp256_ = _2640_ | _2638_;
  assign _2641_ = ~_temp256_;
  assign _2642_ = ~_2641_;
  assign _2643_ = _2642_ ^ _2637_;
  assign _temp257_ = _2643_ ^ _2620_;
  assign _2644_ = ~_temp257_;
  assign _temp258_ = _2534_ | _2532_;
  assign _2645_ = ~_temp258_;
  assign _temp259_ = _2559_ & _2535_;
  assign _temp260_ = _temp259_ | _2645_;
  assign _2646_ = ~_temp260_;
  assign _2647_ = _2646_ ^ _2644_;
  assign _temp261_ = _2553_ | _2539_;
  assign _2648_ = ~_temp261_;
  assign _2649_ = _2558_ & _2554_;
  assign _temp262_ = _2649_ | _2648_;
  assign _2650_ = ~_temp262_;
  assign _2651_ = _2549_ & _2548_;
  assign _2652_ = ~_2551_;
  assign _temp263_ = _2652_ | _2550_;
  assign _2653_ = ~_temp263_;
  assign _temp264_ = _2653_ | _2651_;
  assign _2654_ = ~_temp264_;
  assign _2655_ = b[15] & a[0];
  assign _2656_ = _2655_ ^ _2654_;
  assign _2657_ = _2656_ ^ _2650_;
  assign _temp265_ = _2657_ ^ _2647_;
  assign _2658_ = ~_temp265_;
  assign _temp266_ = _2562_ | _2560_;
  assign _2659_ = ~_temp266_;
  assign _temp267_ = _2568_ & _2563_;
  assign _temp268_ = _temp267_ | _2659_;
  assign _2660_ = ~_temp268_;
  assign _2661_ = _2660_ ^ _2658_;
  assign _2662_ = _2567_ & _2566_;
  assign _2663_ = _2662_ ^ _2661_;
  assign _temp269_ = _2572_ | _2569_;
  assign _2664_ = ~_temp269_;
  assign _2665_ = _2664_ ^ _2663_;
  assign _2666_ = _2574_ & _2573_;
  assign _2667_ = _2666_ ^ _2665_;
  assign _2668_ = _2576_ & _2575_;
  assign _2669_ = _2668_ ^ _2667_;
  assign _2670_ = _2578_ & _2577_;
  assign _temp270_ = _2586_ & _2579_;
  assign _temp271_ = _temp270_ | _2670_;
  assign _2671_ = ~_temp271_;
  assign _temp272_ = _2671_ ^ _2669_;
  assign q[15] = ~_temp272_;
  assign _2672_ = a[16] & b[0];
  assign _2673_ = b[1] & a[15];
  assign _2674_ = _2673_ ^ _2672_;
  assign _2675_ = b[2] & a[14];
  assign _temp273_ = _2675_ ^ _2674_;
  assign _2676_ = ~_temp273_;
  assign _2677_ = _2588_ & _2587_;
  assign _temp274_ = _2590_ & _2589_;
  assign _temp275_ = _temp274_ | _2677_;
  assign _2678_ = ~_temp275_;
  assign _2679_ = _2678_ ^ _2676_;
  assign _2680_ = b[3] & a[13];
  assign _2681_ = b[4] & a[12];
  assign _2682_ = _2681_ ^ _2680_;
  assign _2683_ = b[5] & a[11];
  assign _temp276_ = _2683_ ^ _2682_;
  assign _2684_ = ~_temp276_;
  assign _2685_ = _2684_ ^ _2679_;
  assign _temp277_ = _2593_ | _2591_;
  assign _2686_ = ~_temp277_;
  assign _temp278_ = _2599_ & _2594_;
  assign _temp279_ = _temp278_ | _2686_;
  assign _2687_ = ~_temp279_;
  assign _2688_ = _2687_ ^ _2685_;
  assign _2689_ = _2596_ & _2595_;
  assign _2690_ = _2598_ & _2597_;
  assign _temp280_ = _2690_ | _2689_;
  assign _2691_ = ~_temp280_;
  assign _2692_ = b[6] & a[10];
  assign _2693_ = b[7] & a[9];
  assign _2694_ = _2693_ ^ _2692_;
  assign _2695_ = b[8] & a[8];
  assign _temp281_ = _2695_ ^ _2694_;
  assign _2696_ = ~_temp281_;
  assign _2697_ = _2696_ ^ _2691_;
  assign _2698_ = _2608_ & _2607_;
  assign _2699_ = _2610_ & _2609_;
  assign _2700_ = _2699_ | _2698_;
  assign _2701_ = _2700_ ^ _2697_;
  assign _temp282_ = _2701_ ^ _2688_;
  assign _2702_ = ~_temp282_;
  assign _temp283_ = _2602_ | _2600_;
  assign _2703_ = ~_temp283_;
  assign _temp284_ = _2616_ & _2603_;
  assign _temp285_ = _temp284_ | _2703_;
  assign _2704_ = ~_temp285_;
  assign _2705_ = _2704_ ^ _2702_;
  assign _temp286_ = _2611_ | _2606_;
  assign _2706_ = ~_temp286_;
  assign _2707_ = _2615_ & _2612_;
  assign _temp287_ = _2707_ | _2706_;
  assign _2708_ = ~_temp287_;
  assign _2709_ = b[9] & a[7];
  assign _2710_ = b[10] & a[6];
  assign _2711_ = _2710_ ^ _2709_;
  assign _2712_ = b[11] & a[5];
  assign _temp288_ = _2712_ ^ _2711_;
  assign _2713_ = ~_temp288_;
  assign _2714_ = _2624_ & _2623_;
  assign _temp289_ = _2626_ & _2625_;
  assign _temp290_ = _temp289_ | _2714_;
  assign _2715_ = ~_temp290_;
  assign _2716_ = _2715_ ^ _2713_;
  assign _2717_ = b[12] & a[4];
  assign _2718_ = b[13] & a[3];
  assign _2719_ = _2718_ ^ _2717_;
  assign _2720_ = b[14] & a[2];
  assign _temp291_ = _2720_ ^ _2719_;
  assign _2721_ = ~_temp291_;
  assign _2722_ = _2721_ ^ _2716_;
  assign _temp292_ = _2722_ ^ _2708_;
  assign _2723_ = ~_temp292_;
  assign _temp293_ = _2629_ | _2627_;
  assign _2724_ = ~_temp293_;
  assign _2725_ = ~_2635_;
  assign _2726_ = _2725_ & _2630_;
  assign _temp294_ = _2726_ | _2724_;
  assign _2727_ = ~_temp294_;
  assign _2728_ = _2727_ ^ _2723_;
  assign _temp295_ = _2728_ ^ _2705_;
  assign _2729_ = ~_temp295_;
  assign _temp296_ = _2619_ | _2617_;
  assign _2730_ = ~_temp296_;
  assign _temp297_ = _2643_ & _2620_;
  assign _temp298_ = _temp297_ | _2730_;
  assign _2731_ = ~_temp298_;
  assign _2732_ = _2731_ ^ _2729_;
  assign _temp299_ = _2636_ | _2622_;
  assign _2733_ = ~_temp299_;
  assign _2734_ = _2642_ & _2637_;
  assign _temp300_ = _2734_ | _2733_;
  assign _2735_ = ~_temp300_;
  assign _2736_ = ~_2634_;
  assign _temp301_ = _2632_ & _2631_;
  assign _2737_ = ~_temp301_;
  assign _temp302_ = _2736_ | _2633_;
  assign _temp303_ = _temp302_ & _2737_;
  assign _2738_ = ~_temp303_;
  assign _2739_ = b[15] & a[1];
  assign _2740_ = b[16] & a[0];
  assign _temp304_ = _2740_ ^ _2739_;
  assign _2741_ = ~_temp304_;
  assign _2742_ = _2741_ ^ _2738_;
  assign _2743_ = ~_2655_;
  assign _temp305_ = _2743_ | _2654_;
  assign _2744_ = ~_temp305_;
  assign _2745_ = _2744_ ^ _2742_;
  assign _2746_ = _2745_ ^ _2735_;
  assign _temp306_ = _2746_ ^ _2732_;
  assign _2747_ = ~_temp306_;
  assign _temp307_ = _2646_ | _2644_;
  assign _2748_ = ~_temp307_;
  assign _temp308_ = _2657_ & _2647_;
  assign _temp309_ = _temp308_ | _2748_;
  assign _2749_ = ~_temp309_;
  assign _2750_ = _2749_ ^ _2747_;
  assign _temp310_ = _2656_ | _2650_;
  assign _2751_ = ~_temp310_;
  assign _temp311_ = _2751_ ^ _2750_;
  assign _2752_ = ~_temp311_;
  assign _temp312_ = _2660_ | _2658_;
  assign _2753_ = ~_temp312_;
  assign _temp313_ = _2662_ & _2661_;
  assign _temp314_ = _temp313_ | _2753_;
  assign _2754_ = ~_temp314_;
  assign _2755_ = _2754_ ^ _2752_;
  assign _2756_ = _2664_ & _2663_;
  assign _2757_ = _2756_ ^ _2755_;
  assign _2758_ = _2666_ & _2665_;
  assign _2759_ = _2758_ ^ _2757_;
  assign _2760_ = ~_2759_;
  assign _2761_ = _2669_ & _2579_;
  assign _2762_ = _2761_ & _2585_;
  assign _temp315_ = _2669_ & _2579_;
  assign _2763_ = ~_temp315_;
  assign _2764_ = _2668_ & _2667_;
  assign _temp316_ = _2670_ & _2669_;
  assign _temp317_ = _temp316_ | _2764_;
  assign _2765_ = ~_temp317_;
  assign _temp318_ = _2763_ | _2582_;
  assign _temp319_ = _temp318_ & _2765_;
  assign _2766_ = ~_temp319_;
  assign _temp320_ = _2766_ | _2762_;
  assign _2767_ = ~_temp320_;
  assign q[16] = _2767_ ^ _2760_;
  assign _2768_ = a[17] & b[0];
  assign _2769_ = b[1] & a[16];
  assign _2770_ = _2769_ ^ _2768_;
  assign _2771_ = b[2] & a[15];
  assign _temp321_ = _2771_ ^ _2770_;
  assign _2772_ = ~_temp321_;
  assign _2773_ = _2673_ & _2672_;
  assign _temp322_ = _2675_ & _2674_;
  assign _temp323_ = _temp322_ | _2773_;
  assign _2774_ = ~_temp323_;
  assign _2775_ = _2774_ ^ _2772_;
  assign _2776_ = b[3] & a[14];
  assign _2777_ = b[4] & a[13];
  assign _2778_ = _2777_ ^ _2776_;
  assign _2779_ = b[5] & a[12];
  assign _2780_ = _2779_ ^ _2778_;
  assign _temp324_ = _2780_ ^ _2775_;
  assign _2781_ = ~_temp324_;
  assign _2782_ = ~_2684_;
  assign _temp325_ = _2678_ | _2676_;
  assign _2783_ = ~_temp325_;
  assign _temp326_ = _2782_ & _2679_;
  assign _temp327_ = _temp326_ | _2783_;
  assign _2784_ = ~_temp327_;
  assign _2785_ = _2784_ ^ _2781_;
  assign _2786_ = _2681_ & _2680_;
  assign _2787_ = _2683_ & _2682_;
  assign _temp328_ = _2787_ | _2786_;
  assign _2788_ = ~_temp328_;
  assign _2789_ = b[6] & a[11];
  assign _2790_ = b[7] & a[10];
  assign _2791_ = _2790_ ^ _2789_;
  assign _2792_ = b[8] & a[9];
  assign _temp329_ = _2792_ ^ _2791_;
  assign _2793_ = ~_temp329_;
  assign _2794_ = _2793_ ^ _2788_;
  assign _2795_ = _2693_ & _2692_;
  assign _2796_ = _2695_ & _2694_;
  assign _2797_ = _2796_ | _2795_;
  assign _2798_ = _2797_ ^ _2794_;
  assign _temp330_ = _2798_ ^ _2785_;
  assign _2799_ = ~_temp330_;
  assign _temp331_ = _2687_ | _2685_;
  assign _2800_ = ~_temp331_;
  assign _temp332_ = _2701_ & _2688_;
  assign _temp333_ = _temp332_ | _2800_;
  assign _2801_ = ~_temp333_;
  assign _2802_ = _2801_ ^ _2799_;
  assign _temp334_ = _2696_ | _2691_;
  assign _2803_ = ~_temp334_;
  assign _2804_ = _2700_ & _2697_;
  assign _temp335_ = _2804_ | _2803_;
  assign _2805_ = ~_temp335_;
  assign _2806_ = b[9] & a[8];
  assign _2807_ = b[10] & a[7];
  assign _2808_ = _2807_ ^ _2806_;
  assign _2809_ = b[11] & a[6];
  assign _temp336_ = _2809_ ^ _2808_;
  assign _2810_ = ~_temp336_;
  assign _2811_ = _2710_ & _2709_;
  assign _temp337_ = _2712_ & _2711_;
  assign _temp338_ = _temp337_ | _2811_;
  assign _2812_ = ~_temp338_;
  assign _2813_ = _2812_ ^ _2810_;
  assign _2814_ = b[12] & a[5];
  assign _2815_ = b[13] & a[4];
  assign _2816_ = _2815_ ^ _2814_;
  assign _2817_ = b[14] & a[3];
  assign _temp339_ = _2817_ ^ _2816_;
  assign _2818_ = ~_temp339_;
  assign _2819_ = _2818_ ^ _2813_;
  assign _temp340_ = _2819_ ^ _2805_;
  assign _2820_ = ~_temp340_;
  assign _temp341_ = _2715_ | _2713_;
  assign _2821_ = ~_temp341_;
  assign _2822_ = ~_2721_;
  assign _2823_ = _2822_ & _2716_;
  assign _temp342_ = _2823_ | _2821_;
  assign _2824_ = ~_temp342_;
  assign _2825_ = _2824_ ^ _2820_;
  assign _temp343_ = _2825_ ^ _2802_;
  assign _2826_ = ~_temp343_;
  assign _temp344_ = _2704_ | _2702_;
  assign _2827_ = ~_temp344_;
  assign _temp345_ = _2728_ & _2705_;
  assign _temp346_ = _temp345_ | _2827_;
  assign _2828_ = ~_temp346_;
  assign _2829_ = _2828_ ^ _2826_;
  assign _2830_ = _2722_ ^ _2708_;
  assign _2831_ = ~_2727_;
  assign _temp347_ = _2722_ | _2708_;
  assign _2832_ = ~_temp347_;
  assign _temp348_ = _2831_ & _2830_;
  assign _temp349_ = _temp348_ | _2832_;
  assign _2833_ = ~_temp349_;
  assign _2834_ = _2718_ & _2717_;
  assign _2835_ = _2720_ & _2719_;
  assign _temp350_ = _2835_ | _2834_;
  assign _2836_ = ~_temp350_;
  assign _2837_ = b[15] & a[2];
  assign _2838_ = b[16] & a[1];
  assign _2839_ = _2838_ ^ _2837_;
  assign _2840_ = b[17] & a[0];
  assign _temp351_ = _2840_ ^ _2839_;
  assign _2841_ = ~_temp351_;
  assign _2842_ = _2841_ ^ _2836_;
  assign _2843_ = _2740_ & _2739_;
  assign _temp352_ = _2843_ ^ _2842_;
  assign _2844_ = ~_temp352_;
  assign _2845_ = ~_2741_;
  assign _2846_ = _2845_ & _2738_;
  assign _2847_ = _2846_ ^ _2844_;
  assign _2848_ = _2847_ ^ _2833_;
  assign _2849_ = ~_2742_;
  assign _2850_ = _2744_ & _2849_;
  assign _2851_ = _2850_ ^ _2848_;
  assign _temp353_ = _2851_ ^ _2829_;
  assign _2852_ = ~_temp353_;
  assign _temp354_ = _2731_ | _2729_;
  assign _2853_ = ~_temp354_;
  assign _temp355_ = _2746_ & _2732_;
  assign _temp356_ = _temp355_ | _2853_;
  assign _2854_ = ~_temp356_;
  assign _2855_ = _2854_ ^ _2852_;
  assign _temp357_ = _2745_ | _2735_;
  assign _2856_ = ~_temp357_;
  assign _temp358_ = _2856_ ^ _2855_;
  assign _2857_ = ~_temp358_;
  assign _temp359_ = _2749_ | _2747_;
  assign _2858_ = ~_temp359_;
  assign _temp360_ = _2751_ & _2750_;
  assign _temp361_ = _temp360_ | _2858_;
  assign _2859_ = ~_temp361_;
  assign _2860_ = _2859_ ^ _2857_;
  assign _temp362_ = _2754_ | _2752_;
  assign _2861_ = ~_temp362_;
  assign _2862_ = _2861_ ^ _2860_;
  assign _2863_ = _2756_ & _2755_;
  assign _2864_ = _2863_ ^ _2862_;
  assign _2865_ = _2758_ & _2757_;
  assign _2866_ = ~_2865_;
  assign _temp363_ = _2767_ | _2760_;
  assign _temp364_ = _temp363_ & _2866_;
  assign _2867_ = ~_temp364_;
  assign q[17] = _2867_ ^ _2864_;
  assign _2868_ = a[18] & b[0];
  assign _2869_ = b[1] & a[17];
  assign _2870_ = _2869_ ^ _2868_;
  assign _2871_ = b[2] & a[16];
  assign _temp365_ = _2871_ ^ _2870_;
  assign _2872_ = ~_temp365_;
  assign _2873_ = _2769_ & _2768_;
  assign _temp366_ = _2771_ & _2770_;
  assign _temp367_ = _temp366_ | _2873_;
  assign _2875_ = ~_temp367_;
  assign _2876_ = _2875_ ^ _2872_;
  assign _2877_ = b[3] & a[15];
  assign _2878_ = b[4] & a[14];
  assign _2879_ = _2878_ ^ _2877_;
  assign _2880_ = b[5] & a[13];
  assign _2881_ = _2880_ ^ _2879_;
  assign _temp368_ = _2881_ ^ _2876_;
  assign _2882_ = ~_temp368_;
  assign _temp369_ = _2774_ | _2772_;
  assign _2883_ = ~_temp369_;
  assign _temp370_ = _2780_ & _2775_;
  assign _temp371_ = _temp370_ | _2883_;
  assign _2884_ = ~_temp371_;
  assign _2886_ = _2884_ ^ _2882_;
  assign _2887_ = _2777_ & _2776_;
  assign _2888_ = _2779_ & _2778_;
  assign _temp372_ = _2888_ | _2887_;
  assign _2889_ = ~_temp372_;
  assign _2890_ = b[6] & a[12];
  assign _2891_ = b[7] & a[11];
  assign _2892_ = _2891_ ^ _2890_;
  assign _2893_ = b[8] & a[10];
  assign _temp373_ = _2893_ ^ _2892_;
  assign _2894_ = ~_temp373_;
  assign _temp374_ = _2894_ ^ _2889_;
  assign _2895_ = ~_temp374_;
  assign _2896_ = _2790_ & _2789_;
  assign _2897_ = _2792_ & _2791_;
  assign _temp375_ = _2897_ | _2896_;
  assign _2898_ = ~_temp375_;
  assign _2899_ = _2898_ ^ _2895_;
  assign _temp376_ = _2899_ ^ _2886_;
  assign _2900_ = ~_temp376_;
  assign _temp377_ = _2784_ | _2781_;
  assign _2901_ = ~_temp377_;
  assign _temp378_ = _2798_ & _2785_;
  assign _temp379_ = _temp378_ | _2901_;
  assign _2902_ = ~_temp379_;
  assign _2903_ = _2902_ ^ _2900_;
  assign _temp380_ = _2793_ | _2788_;
  assign _2904_ = ~_temp380_;
  assign _2905_ = _2797_ & _2794_;
  assign _temp381_ = _2905_ | _2904_;
  assign _0000_ = ~_temp381_;
  assign _0001_ = b[9] & a[9];
  assign _0002_ = b[10] & a[8];
  assign _0003_ = _0002_ ^ _0001_;
  assign _0004_ = b[11] & a[7];
  assign _temp382_ = _0004_ ^ _0003_;
  assign _0005_ = ~_temp382_;
  assign _0006_ = _2807_ & _2806_;
  assign _temp383_ = _2809_ & _2808_;
  assign _temp384_ = _temp383_ | _0006_;
  assign _0007_ = ~_temp384_;
  assign _0008_ = _0007_ ^ _0005_;
  assign _0009_ = b[12] & a[6];
  assign _0011_ = b[13] & a[5];
  assign _0012_ = _0011_ ^ _0009_;
  assign _0013_ = b[14] & a[4];
  assign _temp385_ = _0013_ ^ _0012_;
  assign _0014_ = ~_temp385_;
  assign _0015_ = _0014_ ^ _0008_;
  assign _temp386_ = _0015_ ^ _0000_;
  assign _0016_ = ~_temp386_;
  assign _temp387_ = _2812_ | _2810_;
  assign _0017_ = ~_temp387_;
  assign _0018_ = ~_2818_;
  assign _0019_ = _0018_ & _2813_;
  assign _temp388_ = _0019_ | _0017_;
  assign _0020_ = ~_temp388_;
  assign _0022_ = _0020_ ^ _0016_;
  assign _temp389_ = _0022_ ^ _2903_;
  assign _0023_ = ~_temp389_;
  assign _temp390_ = _2801_ | _2799_;
  assign _0024_ = ~_temp390_;
  assign _temp391_ = _2825_ & _2802_;
  assign _temp392_ = _temp391_ | _0024_;
  assign _0025_ = ~_temp392_;
  assign _0026_ = _0025_ ^ _0023_;
  assign _0027_ = _2819_ ^ _2805_;
  assign _0028_ = ~_2824_;
  assign _temp393_ = _2819_ | _2805_;
  assign _0029_ = ~_temp393_;
  assign _temp394_ = _0028_ & _0027_;
  assign _temp395_ = _temp394_ | _0029_;
  assign _0030_ = ~_temp395_;
  assign _0031_ = _2815_ & _2814_;
  assign _0033_ = _2817_ & _2816_;
  assign _temp396_ = _0033_ | _0031_;
  assign _0034_ = ~_temp396_;
  assign _0035_ = b[15] & a[3];
  assign _0036_ = b[16] & a[2];
  assign _0037_ = _0036_ ^ _0035_;
  assign _0038_ = b[17] & a[1];
  assign _temp397_ = _0038_ ^ _0037_;
  assign _0039_ = ~_temp397_;
  assign _0040_ = _0039_ ^ _0034_;
  assign _0041_ = _2838_ & _2837_;
  assign _0042_ = _2840_ & _2839_;
  assign _0044_ = _0042_ | _0041_;
  assign _temp398_ = _0044_ ^ _0040_;
  assign _0045_ = ~_temp398_;
  assign _temp399_ = _2841_ | _2836_;
  assign _0046_ = ~_temp399_;
  assign _temp400_ = _2843_ & _2842_;
  assign _temp401_ = _temp400_ | _0046_;
  assign _0047_ = ~_temp401_;
  assign _0048_ = _0047_ ^ _0045_;
  assign _0049_ = b[18] & a[0];
  assign _temp402_ = _0049_ ^ _0048_;
  assign _0050_ = ~_temp402_;
  assign _0051_ = _0050_ ^ _0030_;
  assign _0052_ = ~_2846_;
  assign _temp403_ = _0052_ | _2844_;
  assign _0053_ = ~_temp403_;
  assign _0055_ = _0053_ ^ _0051_;
  assign _temp404_ = _0055_ ^ _0026_;
  assign _0056_ = ~_temp404_;
  assign _temp405_ = _2828_ | _2826_;
  assign _0057_ = ~_temp405_;
  assign _temp406_ = _2851_ & _2829_;
  assign _temp407_ = _temp406_ | _0057_;
  assign _0058_ = ~_temp407_;
  assign _0059_ = _0058_ ^ _0056_;
  assign _temp408_ = _2847_ | _2833_;
  assign _0060_ = ~_temp408_;
  assign _0061_ = _2850_ & _2848_;
  assign _0062_ = _0061_ | _0060_;
  assign _temp409_ = _0062_ ^ _0059_;
  assign _0063_ = ~_temp409_;
  assign _temp410_ = _2854_ | _2852_;
  assign _0064_ = ~_temp410_;
  assign _temp411_ = _2856_ & _2855_;
  assign _temp412_ = _temp411_ | _0064_;
  assign _0066_ = ~_temp412_;
  assign _0067_ = _0066_ ^ _0063_;
  assign _temp413_ = _2859_ | _2857_;
  assign _0068_ = ~_temp413_;
  assign _0069_ = _0068_ ^ _0067_;
  assign _0070_ = _2861_ & _2860_;
  assign _0071_ = _0070_ ^ _0069_;
  assign _0072_ = _2863_ & _2862_;
  assign _temp414_ = _2865_ & _2864_;
  assign _temp415_ = _temp414_ | _0072_;
  assign _0073_ = ~_temp415_;
  assign _temp416_ = _2864_ & _2759_;
  assign _0074_ = ~_temp416_;
  assign _temp417_ = _0074_ | _2767_;
  assign _temp418_ = _temp417_ & _0073_;
  assign _0075_ = ~_temp418_;
  assign q[18] = _0075_ ^ _0071_;
  assign _0077_ = a[19] & b[0];
  assign _0078_ = b[1] & a[18];
  assign _0079_ = _0078_ ^ _0077_;
  assign _0080_ = b[2] & a[17];
  assign _temp419_ = _0080_ ^ _0079_;
  assign _0081_ = ~_temp419_;
  assign _0082_ = _2869_ & _2868_;
  assign _temp420_ = _2871_ & _2870_;
  assign _temp421_ = _temp420_ | _0082_;
  assign _0083_ = ~_temp421_;
  assign _0084_ = _0083_ ^ _0081_;
  assign _0085_ = b[3] & a[16];
  assign _0086_ = b[4] & a[15];
  assign _0087_ = _0086_ ^ _0085_;
  assign _0088_ = b[5] & a[14];
  assign _0089_ = _0088_ ^ _0087_;
  assign _temp422_ = _0089_ ^ _0084_;
  assign _0090_ = ~_temp422_;
  assign _temp423_ = _2875_ | _2872_;
  assign _0091_ = ~_temp423_;
  assign _temp424_ = _2881_ & _2876_;
  assign _temp425_ = _temp424_ | _0091_;
  assign _0092_ = ~_temp425_;
  assign _0093_ = _0092_ ^ _0090_;
  assign _0094_ = _2878_ & _2877_;
  assign _0095_ = _2880_ & _2879_;
  assign _temp426_ = _0095_ | _0094_;
  assign _0097_ = ~_temp426_;
  assign _0098_ = b[6] & a[13];
  assign _0099_ = b[7] & a[12];
  assign _0100_ = _0099_ ^ _0098_;
  assign _0101_ = b[8] & a[11];
  assign _temp427_ = _0101_ ^ _0100_;
  assign _0102_ = ~_temp427_;
  assign _temp428_ = _0102_ ^ _0097_;
  assign _0103_ = ~_temp428_;
  assign _0104_ = _2891_ & _2890_;
  assign _0105_ = _2893_ & _2892_;
  assign _temp429_ = _0105_ | _0104_;
  assign _0106_ = ~_temp429_;
  assign _0108_ = _0106_ ^ _0103_;
  assign _temp430_ = _0108_ ^ _0093_;
  assign _0109_ = ~_temp430_;
  assign _temp431_ = _2884_ | _2882_;
  assign _0110_ = ~_temp431_;
  assign _temp432_ = _2899_ & _2886_;
  assign _temp433_ = _temp432_ | _0110_;
  assign _0111_ = ~_temp433_;
  assign _0112_ = _0111_ ^ _0109_;
  assign _0113_ = _2894_ ^ _2889_;
  assign _0114_ = _2897_ | _2896_;
  assign _temp434_ = _2894_ | _2889_;
  assign _0115_ = ~_temp434_;
  assign _temp435_ = _0114_ & _0113_;
  assign _temp436_ = _temp435_ | _0115_;
  assign _0116_ = ~_temp436_;
  assign _0117_ = b[9] & a[10];
  assign _0119_ = b[10] & a[9];
  assign _0120_ = _0119_ ^ _0117_;
  assign _0121_ = b[11] & a[8];
  assign _temp437_ = _0121_ ^ _0120_;
  assign _0122_ = ~_temp437_;
  assign _0123_ = _0002_ & _0001_;
  assign _temp438_ = _0004_ & _0003_;
  assign _temp439_ = _temp438_ | _0123_;
  assign _0124_ = ~_temp439_;
  assign _0125_ = _0124_ ^ _0122_;
  assign _0126_ = b[12] & a[7];
  assign _0127_ = b[13] & a[6];
  assign _0128_ = _0127_ ^ _0126_;
  assign _0130_ = b[14] & a[5];
  assign _temp440_ = _0130_ ^ _0128_;
  assign _0131_ = ~_temp440_;
  assign _0132_ = _0131_ ^ _0125_;
  assign _temp441_ = _0132_ ^ _0116_;
  assign _0133_ = ~_temp441_;
  assign _temp442_ = _0007_ | _0005_;
  assign _0134_ = ~_temp442_;
  assign _0135_ = ~_0014_;
  assign _0136_ = _0135_ & _0008_;
  assign _temp443_ = _0136_ | _0134_;
  assign _0137_ = ~_temp443_;
  assign _0138_ = _0137_ ^ _0133_;
  assign _temp444_ = _0138_ ^ _0112_;
  assign _0139_ = ~_temp444_;
  assign _temp445_ = _2902_ | _2900_;
  assign _0141_ = ~_temp445_;
  assign _temp446_ = _0022_ & _2903_;
  assign _temp447_ = _temp446_ | _0141_;
  assign _0142_ = ~_temp447_;
  assign _0143_ = _0142_ ^ _0139_;
  assign _0144_ = _0015_ ^ _0000_;
  assign _0145_ = ~_0020_;
  assign _temp448_ = _0015_ | _0000_;
  assign _0146_ = ~_temp448_;
  assign _temp449_ = _0145_ & _0144_;
  assign _temp450_ = _temp449_ | _0146_;
  assign _0147_ = ~_temp450_;
  assign _0148_ = _0011_ & _0009_;
  assign _temp451_ = _0013_ & _0012_;
  assign _temp452_ = _temp451_ | _0148_;
  assign _0149_ = ~_temp452_;
  assign _0150_ = b[15] & a[4];
  assign _0152_ = b[16] & a[3];
  assign _0153_ = _0152_ ^ _0150_;
  assign _0154_ = b[17] & a[2];
  assign _temp453_ = _0154_ ^ _0153_;
  assign _0155_ = ~_temp453_;
  assign _0156_ = _0155_ ^ _0149_;
  assign _0157_ = _0036_ & _0035_;
  assign _0158_ = _0038_ & _0037_;
  assign _0159_ = _0158_ | _0157_;
  assign _temp454_ = _0159_ ^ _0156_;
  assign _0160_ = ~_temp454_;
  assign _temp455_ = _0039_ | _0034_;
  assign _0161_ = ~_temp455_;
  assign _temp456_ = _0044_ & _0040_;
  assign _temp457_ = _temp456_ | _0161_;
  assign _0163_ = ~_temp457_;
  assign _0164_ = _0163_ ^ _0160_;
  assign _0165_ = b[18] & a[1];
  assign _0166_ = b[19] & a[0];
  assign _temp458_ = _0166_ ^ _0165_;
  assign _0167_ = ~_temp458_;
  assign _0168_ = _0167_ ^ _0164_;
  assign _0169_ = _0168_ ^ _0147_;
  assign _temp459_ = _0047_ | _0045_;
  assign _0170_ = ~_temp459_;
  assign _0171_ = _0049_ & _0048_;
  assign _temp460_ = _0171_ | _0170_;
  assign _0172_ = ~_temp460_;
  assign _0174_ = ~_0172_;
  assign _0175_ = _0174_ ^ _0169_;
  assign _temp461_ = _0175_ ^ _0143_;
  assign _0176_ = ~_temp461_;
  assign _temp462_ = _0025_ | _0023_;
  assign _0177_ = ~_temp462_;
  assign _temp463_ = _0055_ & _0026_;
  assign _temp464_ = _temp463_ | _0177_;
  assign _0178_ = ~_temp464_;
  assign _0179_ = _0178_ ^ _0176_;
  assign _temp465_ = _0050_ | _0030_;
  assign _0180_ = ~_temp465_;
  assign _0181_ = _0053_ & _0051_;
  assign _0182_ = _0181_ | _0180_;
  assign _temp466_ = _0182_ ^ _0179_;
  assign _0183_ = ~_temp466_;
  assign _temp467_ = _0058_ | _0056_;
  assign _0185_ = ~_temp467_;
  assign _temp468_ = _0062_ & _0059_;
  assign _temp469_ = _temp468_ | _0185_;
  assign _0186_ = ~_temp469_;
  assign _0187_ = _0186_ ^ _0183_;
  assign _temp470_ = _0066_ | _0063_;
  assign _0188_ = ~_temp470_;
  assign _0189_ = _0188_ ^ _0187_;
  assign _0190_ = _0068_ & _0067_;
  assign _0191_ = _0190_ ^ _0189_;
  assign _0192_ = _0070_ & _0069_;
  assign _temp471_ = _0075_ & _0071_;
  assign _temp472_ = _temp471_ | _0192_;
  assign _0193_ = ~_temp472_;
  assign _temp473_ = _0193_ ^ _0191_;
  assign q[19] = ~_temp473_;
  assign _0195_ = a[20] & b[0];
  assign _0196_ = b[1] & a[19];
  assign _0197_ = _0196_ ^ _0195_;
  assign _0198_ = b[2] & a[18];
  assign _temp474_ = _0198_ ^ _0197_;
  assign _0199_ = ~_temp474_;
  assign _0200_ = _0078_ & _0077_;
  assign _temp475_ = _0080_ & _0079_;
  assign _temp476_ = _temp475_ | _0200_;
  assign _0201_ = ~_temp476_;
  assign _0202_ = _0201_ ^ _0199_;
  assign _0203_ = b[3] & a[17];
  assign _0204_ = b[4] & a[16];
  assign _0206_ = _0204_ ^ _0203_;
  assign _0207_ = b[5] & a[15];
  assign _0208_ = _0207_ ^ _0206_;
  assign _temp477_ = _0208_ ^ _0202_;
  assign _0209_ = ~_temp477_;
  assign _temp478_ = _0083_ | _0081_;
  assign _0210_ = ~_temp478_;
  assign _temp479_ = _0089_ & _0084_;
  assign _temp480_ = _temp479_ | _0210_;
  assign _0211_ = ~_temp480_;
  assign _0212_ = _0211_ ^ _0209_;
  assign _0213_ = _0086_ & _0085_;
  assign _0214_ = _0088_ & _0087_;
  assign _temp481_ = _0214_ | _0213_;
  assign _0215_ = ~_temp481_;
  assign _0217_ = b[6] & a[14];
  assign _0218_ = b[7] & a[13];
  assign _0219_ = _0218_ ^ _0217_;
  assign _0220_ = b[8] & a[12];
  assign _temp482_ = _0220_ ^ _0219_;
  assign _0221_ = ~_temp482_;
  assign _temp483_ = _0221_ ^ _0215_;
  assign _0222_ = ~_temp483_;
  assign _0223_ = _0099_ & _0098_;
  assign _0224_ = _0101_ & _0100_;
  assign _temp484_ = _0224_ | _0223_;
  assign _0225_ = ~_temp484_;
  assign _0226_ = _0225_ ^ _0222_;
  assign _temp485_ = _0226_ ^ _0212_;
  assign _0227_ = ~_temp485_;
  assign _temp486_ = _0092_ | _0090_;
  assign _0228_ = ~_temp486_;
  assign _temp487_ = _0108_ & _0093_;
  assign _temp488_ = _temp487_ | _0228_;
  assign _0229_ = ~_temp488_;
  assign _0230_ = _0229_ ^ _0227_;
  assign _0231_ = _0102_ ^ _0097_;
  assign _0232_ = _0105_ | _0104_;
  assign _temp489_ = _0102_ | _0097_;
  assign _0233_ = ~_temp489_;
  assign _temp490_ = _0232_ & _0231_;
  assign _temp491_ = _temp490_ | _0233_;
  assign _0234_ = ~_temp491_;
  assign _0235_ = b[9] & a[11];
  assign _0236_ = b[10] & a[10];
  assign _0238_ = _0236_ ^ _0235_;
  assign _0239_ = b[11] & a[9];
  assign _temp492_ = _0239_ ^ _0238_;
  assign _0240_ = ~_temp492_;
  assign _0241_ = _0119_ & _0117_;
  assign _temp493_ = _0121_ & _0120_;
  assign _temp494_ = _temp493_ | _0241_;
  assign _0242_ = ~_temp494_;
  assign _0243_ = _0242_ ^ _0240_;
  assign _0244_ = b[12] & a[8];
  assign _0245_ = b[13] & a[7];
  assign _0246_ = _0245_ ^ _0244_;
  assign _0247_ = b[14] & a[6];
  assign _temp495_ = _0247_ ^ _0246_;
  assign _0249_ = ~_temp495_;
  assign _0250_ = _0249_ ^ _0243_;
  assign _temp496_ = _0250_ ^ _0234_;
  assign _0251_ = ~_temp496_;
  assign _temp497_ = _0124_ | _0122_;
  assign _0252_ = ~_temp497_;
  assign _0253_ = ~_0131_;
  assign _0254_ = _0253_ & _0125_;
  assign _temp498_ = _0254_ | _0252_;
  assign _0255_ = ~_temp498_;
  assign _0256_ = _0255_ ^ _0251_;
  assign _temp499_ = _0256_ ^ _0230_;
  assign _0257_ = ~_temp499_;
  assign _temp500_ = _0111_ | _0109_;
  assign _0258_ = ~_temp500_;
  assign _temp501_ = _0138_ & _0112_;
  assign _temp502_ = _temp501_ | _0258_;
  assign _0260_ = ~_temp502_;
  assign _0261_ = _0260_ ^ _0257_;
  assign _0262_ = _0132_ | _0116_;
  assign _temp503_ = _0137_ | _0133_;
  assign _temp504_ = _temp503_ & _0262_;
  assign _0263_ = ~_temp504_;
  assign _0264_ = _0127_ & _0126_;
  assign _temp505_ = _0130_ & _0128_;
  assign _temp506_ = _temp505_ | _0264_;
  assign _0265_ = ~_temp506_;
  assign _0266_ = b[15] & a[5];
  assign _0267_ = b[16] & a[4];
  assign _0268_ = _0267_ ^ _0266_;
  assign _0269_ = b[17] & a[3];
  assign _temp507_ = _0269_ ^ _0268_;
  assign _0271_ = ~_temp507_;
  assign _0272_ = _0271_ ^ _0265_;
  assign _0273_ = _0152_ & _0150_;
  assign _0274_ = _0154_ & _0153_;
  assign _0275_ = _0274_ | _0273_;
  assign _temp508_ = _0275_ ^ _0272_;
  assign _0276_ = ~_temp508_;
  assign _temp509_ = _0155_ | _0149_;
  assign _0277_ = ~_temp509_;
  assign _temp510_ = _0159_ & _0156_;
  assign _temp511_ = _temp510_ | _0277_;
  assign _0278_ = ~_temp511_;
  assign _0279_ = _0278_ ^ _0276_;
  assign _0280_ = b[18] & a[2];
  assign _0282_ = b[19] & a[1];
  assign _0283_ = _0282_ ^ _0280_;
  assign _0284_ = b[20] & a[0];
  assign _temp512_ = _0284_ ^ _0283_;
  assign _0285_ = ~_temp512_;
  assign _0286_ = _0166_ & _0165_;
  assign _0287_ = _0286_ ^ _0285_;
  assign _0288_ = _0287_ ^ _0279_;
  assign _0289_ = _0288_ ^ _0263_;
  assign _0290_ = ~_0167_;
  assign _temp513_ = _0163_ | _0160_;
  assign _0291_ = ~_temp513_;
  assign _temp514_ = _0290_ & _0164_;
  assign _temp515_ = _temp514_ | _0291_;
  assign _0293_ = ~_temp515_;
  assign _0294_ = _0293_ ^ _0289_;
  assign _temp516_ = _0294_ ^ _0261_;
  assign _0295_ = ~_temp516_;
  assign _temp517_ = _0142_ | _0139_;
  assign _0296_ = ~_temp517_;
  assign _temp518_ = _0175_ & _0143_;
  assign _temp519_ = _temp518_ | _0296_;
  assign _0297_ = ~_temp519_;
  assign _0298_ = _0297_ ^ _0295_;
  assign _temp520_ = _0168_ | _0147_;
  assign _0299_ = ~_temp520_;
  assign _0300_ = _0174_ & _0169_;
  assign _0301_ = _0300_ | _0299_;
  assign _temp521_ = _0301_ ^ _0298_;
  assign _0302_ = ~_temp521_;
  assign _temp522_ = _0178_ | _0176_;
  assign _0304_ = ~_temp522_;
  assign _temp523_ = _0182_ & _0179_;
  assign _temp524_ = _temp523_ | _0304_;
  assign _0305_ = ~_temp524_;
  assign _0306_ = _0305_ ^ _0302_;
  assign _temp525_ = _0186_ | _0183_;
  assign _0307_ = ~_temp525_;
  assign _0308_ = _0307_ ^ _0306_;
  assign _0309_ = _0188_ & _0187_;
  assign _temp526_ = _0309_ ^ _0308_;
  assign _0310_ = ~_temp526_;
  assign _temp527_ = _0191_ & _0071_;
  assign _0311_ = ~_temp527_;
  assign _0312_ = _0190_ & _0189_;
  assign _temp528_ = _0192_ & _0191_;
  assign _temp529_ = _temp528_ | _0312_;
  assign _0313_ = ~_temp529_;
  assign _temp530_ = _0311_ | _0073_;
  assign _temp531_ = _temp530_ & _0313_;
  assign _0315_ = ~_temp531_;
  assign _0316_ = ~_0315_;
  assign _temp532_ = _0311_ | _0074_;
  assign _0317_ = ~_temp532_;
  assign _temp533_ = _2766_ | _2762_;
  assign _temp534_ = _temp533_ & _0317_;
  assign _0318_ = ~_temp534_;
  assign _0319_ = _0318_ & _0316_;
  assign q[20] = _0319_ ^ _0310_;
  assign _0320_ = a[21] & b[0];
  assign _0321_ = b[1] & a[20];
  assign _0322_ = _0321_ ^ _0320_;
  assign _0323_ = b[2] & a[19];
  assign _temp535_ = _0323_ ^ _0322_;
  assign _0325_ = ~_temp535_;
  assign _0326_ = _0196_ & _0195_;
  assign _temp536_ = _0198_ & _0197_;
  assign _temp537_ = _temp536_ | _0326_;
  assign _0327_ = ~_temp537_;
  assign _0328_ = _0327_ ^ _0325_;
  assign _0329_ = b[3] & a[18];
  assign _0330_ = b[4] & a[17];
  assign _0331_ = _0330_ ^ _0329_;
  assign _0332_ = b[5] & a[16];
  assign _0333_ = _0332_ ^ _0331_;
  assign _temp538_ = _0333_ ^ _0328_;
  assign _0334_ = ~_temp538_;
  assign _temp539_ = _0201_ | _0199_;
  assign _0336_ = ~_temp539_;
  assign _temp540_ = _0208_ & _0202_;
  assign _temp541_ = _temp540_ | _0336_;
  assign _0337_ = ~_temp541_;
  assign _0338_ = _0337_ ^ _0334_;
  assign _0339_ = _0204_ & _0203_;
  assign _0340_ = _0207_ & _0206_;
  assign _temp542_ = _0340_ | _0339_;
  assign _0341_ = ~_temp542_;
  assign _0342_ = b[6] & a[15];
  assign _0343_ = b[7] & a[14];
  assign _0344_ = _0343_ ^ _0342_;
  assign _0345_ = b[8] & a[13];
  assign _temp543_ = _0345_ ^ _0344_;
  assign _0347_ = ~_temp543_;
  assign _temp544_ = _0347_ ^ _0341_;
  assign _0348_ = ~_temp544_;
  assign _0349_ = _0218_ & _0217_;
  assign _0350_ = _0220_ & _0219_;
  assign _temp545_ = _0350_ | _0349_;
  assign _0351_ = ~_temp545_;
  assign _0352_ = _0351_ ^ _0348_;
  assign _temp546_ = _0352_ ^ _0338_;
  assign _0353_ = ~_temp546_;
  assign _temp547_ = _0211_ | _0209_;
  assign _0354_ = ~_temp547_;
  assign _temp548_ = _0226_ & _0212_;
  assign _temp549_ = _temp548_ | _0354_;
  assign _0355_ = ~_temp549_;
  assign _0356_ = _0355_ ^ _0353_;
  assign _0358_ = _0221_ ^ _0215_;
  assign _0359_ = _0224_ | _0223_;
  assign _temp550_ = _0221_ | _0215_;
  assign _0360_ = ~_temp550_;
  assign _temp551_ = _0359_ & _0358_;
  assign _temp552_ = _temp551_ | _0360_;
  assign _0361_ = ~_temp552_;
  assign _0362_ = b[9] & a[12];
  assign _0363_ = b[10] & a[11];
  assign _0364_ = _0363_ ^ _0362_;
  assign _0365_ = b[11] & a[10];
  assign _temp553_ = _0365_ ^ _0364_;
  assign _0366_ = ~_temp553_;
  assign _0367_ = _0236_ & _0235_;
  assign _temp554_ = _0239_ & _0238_;
  assign _temp555_ = _temp554_ | _0367_;
  assign _0369_ = ~_temp555_;
  assign _0370_ = _0369_ ^ _0366_;
  assign _0371_ = b[12] & a[9];
  assign _0372_ = b[13] & a[8];
  assign _0373_ = _0372_ ^ _0371_;
  assign _0374_ = b[14] & a[7];
  assign _temp556_ = _0374_ ^ _0373_;
  assign _0375_ = ~_temp556_;
  assign _0376_ = _0375_ ^ _0370_;
  assign _temp557_ = _0376_ ^ _0361_;
  assign _0377_ = ~_temp557_;
  assign _temp558_ = _0242_ | _0240_;
  assign _0378_ = ~_temp558_;
  assign _0380_ = ~_0249_;
  assign _0381_ = _0380_ & _0243_;
  assign _temp559_ = _0381_ | _0378_;
  assign _0382_ = ~_temp559_;
  assign _0383_ = _0382_ ^ _0377_;
  assign _temp560_ = _0383_ ^ _0356_;
  assign _0384_ = ~_temp560_;
  assign _temp561_ = _0229_ | _0227_;
  assign _0385_ = ~_temp561_;
  assign _temp562_ = _0256_ & _0230_;
  assign _temp563_ = _temp562_ | _0385_;
  assign _0386_ = ~_temp563_;
  assign _0387_ = _0386_ ^ _0384_;
  assign _0388_ = _0250_ ^ _0234_;
  assign _0389_ = _0254_ | _0252_;
  assign _temp564_ = _0250_ | _0234_;
  assign _0391_ = ~_temp564_;
  assign _temp565_ = _0389_ & _0388_;
  assign _temp566_ = _temp565_ | _0391_;
  assign _0392_ = ~_temp566_;
  assign _0393_ = _0245_ & _0244_;
  assign _temp567_ = _0247_ & _0246_;
  assign _temp568_ = _temp567_ | _0393_;
  assign _0394_ = ~_temp568_;
  assign _0395_ = b[15] & a[6];
  assign _0396_ = b[16] & a[5];
  assign _0397_ = _0396_ ^ _0395_;
  assign _0398_ = b[17] & a[4];
  assign _temp569_ = _0398_ ^ _0397_;
  assign _0399_ = ~_temp569_;
  assign _0400_ = _0399_ ^ _0394_;
  assign _0402_ = _0267_ & _0266_;
  assign _0403_ = _0269_ & _0268_;
  assign _0404_ = _0403_ | _0402_;
  assign _temp570_ = _0404_ ^ _0400_;
  assign _0405_ = ~_temp570_;
  assign _temp571_ = _0271_ | _0265_;
  assign _0406_ = ~_temp571_;
  assign _temp572_ = _0275_ & _0272_;
  assign _temp573_ = _temp572_ | _0406_;
  assign _0407_ = ~_temp573_;
  assign _0408_ = _0407_ ^ _0405_;
  assign _0409_ = b[18] & a[3];
  assign _0410_ = b[19] & a[2];
  assign _0411_ = _0410_ ^ _0409_;
  assign _0412_ = b[20] & a[1];
  assign _temp574_ = _0412_ ^ _0411_;
  assign _0413_ = ~_temp574_;
  assign _0414_ = _0282_ & _0280_;
  assign _temp575_ = _0284_ & _0283_;
  assign _temp576_ = _temp575_ | _0414_;
  assign _0415_ = ~_temp576_;
  assign _temp577_ = _0415_ ^ _0413_;
  assign _0416_ = ~_temp577_;
  assign _0417_ = b[21] & a[0];
  assign _0418_ = _0417_ ^ _0416_;
  assign _0419_ = _0418_ ^ _0408_;
  assign _0420_ = _0419_ ^ _0392_;
  assign _temp578_ = _0278_ | _0276_;
  assign _0421_ = ~_temp578_;
  assign _0423_ = ~_0287_;
  assign _0424_ = _0423_ & _0279_;
  assign _0425_ = _0424_ | _0421_;
  assign _0426_ = _0425_ ^ _0420_;
  assign _temp579_ = _0426_ ^ _0387_;
  assign _0427_ = ~_temp579_;
  assign _temp580_ = _0260_ | _0257_;
  assign _0428_ = ~_temp580_;
  assign _temp581_ = _0294_ & _0261_;
  assign _temp582_ = _temp581_ | _0428_;
  assign _0429_ = ~_temp582_;
  assign _0430_ = _0429_ ^ _0427_;
  assign _0431_ = _0137_ | _0133_;
  assign _temp583_ = _0431_ & _0262_;
  assign _temp584_ = _temp583_ | _0288_;
  assign _0432_ = ~_temp584_;
  assign _temp585_ = _0293_ | _0289_;
  assign _0434_ = ~_temp585_;
  assign _0435_ = _0434_ | _0432_;
  assign _0436_ = ~_0286_;
  assign _temp586_ = _0436_ | _0285_;
  assign _0437_ = ~_temp586_;
  assign _0438_ = _0437_ ^ _0435_;
  assign _temp587_ = _0438_ ^ _0430_;
  assign _0439_ = ~_temp587_;
  assign _temp588_ = _0297_ | _0295_;
  assign _0440_ = ~_temp588_;
  assign _temp589_ = _0301_ & _0298_;
  assign _temp590_ = _temp589_ | _0440_;
  assign _0441_ = ~_temp590_;
  assign _0442_ = _0441_ ^ _0439_;
  assign _temp591_ = _0305_ | _0302_;
  assign _0443_ = ~_temp591_;
  assign _0445_ = _0443_ ^ _0442_;
  assign _0446_ = _0307_ & _0306_;
  assign _0447_ = _0446_ ^ _0445_;
  assign _0448_ = _0309_ & _0308_;
  assign _temp592_ = _0319_ | _0310_;
  assign _0449_ = ~_temp592_;
  assign _0450_ = _0449_ | _0448_;
  assign q[21] = _0450_ ^ _0447_;
  assign _0451_ = a[22] & b[0];
  assign _0452_ = b[1] & a[21];
  assign _0453_ = _0452_ ^ _0451_;
  assign _0455_ = b[2] & a[20];
  assign _temp593_ = _0455_ ^ _0453_;
  assign _0456_ = ~_temp593_;
  assign _0457_ = _0321_ & _0320_;
  assign _temp594_ = _0323_ & _0322_;
  assign _temp595_ = _temp594_ | _0457_;
  assign _0458_ = ~_temp595_;
  assign _0459_ = _0458_ ^ _0456_;
  assign _0460_ = b[3] & a[19];
  assign _0461_ = b[4] & a[18];
  assign _0462_ = _0461_ ^ _0460_;
  assign _0463_ = b[5] & a[17];
  assign _0464_ = _0463_ ^ _0462_;
  assign _temp596_ = _0464_ ^ _0459_;
  assign _0466_ = ~_temp596_;
  assign _temp597_ = _0327_ | _0325_;
  assign _0467_ = ~_temp597_;
  assign _temp598_ = _0333_ & _0328_;
  assign _temp599_ = _temp598_ | _0467_;
  assign _0468_ = ~_temp599_;
  assign _0469_ = _0468_ ^ _0466_;
  assign _0470_ = _0330_ & _0329_;
  assign _0471_ = _0332_ & _0331_;
  assign _temp600_ = _0471_ | _0470_;
  assign _0472_ = ~_temp600_;
  assign _0473_ = b[6] & a[16];
  assign _0474_ = b[7] & a[15];
  assign _0475_ = _0474_ ^ _0473_;
  assign _0477_ = b[8] & a[14];
  assign _temp601_ = _0477_ ^ _0475_;
  assign _0478_ = ~_temp601_;
  assign _0479_ = _0478_ ^ _0472_;
  assign _0480_ = _0343_ & _0342_;
  assign _0481_ = _0345_ & _0344_;
  assign _0482_ = _0481_ | _0480_;
  assign _0483_ = _0482_ ^ _0479_;
  assign _temp602_ = _0483_ ^ _0469_;
  assign _0484_ = ~_temp602_;
  assign _temp603_ = _0337_ | _0334_;
  assign _0485_ = ~_temp603_;
  assign _temp604_ = _0352_ & _0338_;
  assign _temp605_ = _temp604_ | _0485_;
  assign _0486_ = ~_temp605_;
  assign _0488_ = _0486_ ^ _0484_;
  assign _0489_ = _0347_ ^ _0341_;
  assign _0490_ = _0350_ | _0349_;
  assign _temp606_ = _0347_ | _0341_;
  assign _0491_ = ~_temp606_;
  assign _temp607_ = _0490_ & _0489_;
  assign _temp608_ = _temp607_ | _0491_;
  assign _0492_ = ~_temp608_;
  assign _0493_ = b[9] & a[13];
  assign _0494_ = b[10] & a[12];
  assign _0495_ = _0494_ ^ _0493_;
  assign _0496_ = b[11] & a[11];
  assign _temp609_ = _0496_ ^ _0495_;
  assign _0497_ = ~_temp609_;
  assign _0499_ = _0363_ & _0362_;
  assign _temp610_ = _0365_ & _0364_;
  assign _temp611_ = _temp610_ | _0499_;
  assign _0500_ = ~_temp611_;
  assign _0501_ = _0500_ ^ _0497_;
  assign _0502_ = b[12] & a[10];
  assign _0503_ = b[13] & a[9];
  assign _0504_ = _0503_ ^ _0502_;
  assign _0505_ = b[14] & a[8];
  assign _temp612_ = _0505_ ^ _0504_;
  assign _0506_ = ~_temp612_;
  assign _0507_ = _0506_ ^ _0501_;
  assign _0508_ = _0507_ ^ _0492_;
  assign _temp613_ = _0369_ | _0366_;
  assign _0510_ = ~_temp613_;
  assign _0511_ = ~_0375_;
  assign _0512_ = _0511_ & _0370_;
  assign _0513_ = _0512_ | _0510_;
  assign _0514_ = _0513_ ^ _0508_;
  assign _temp614_ = _0514_ ^ _0488_;
  assign _0515_ = ~_temp614_;
  assign _temp615_ = _0355_ | _0353_;
  assign _0516_ = ~_temp615_;
  assign _temp616_ = _0383_ & _0356_;
  assign _temp617_ = _temp616_ | _0516_;
  assign _0517_ = ~_temp617_;
  assign _0518_ = _0517_ ^ _0515_;
  assign _0519_ = _0376_ ^ _0361_;
  assign _0521_ = _0381_ | _0378_;
  assign _temp618_ = _0376_ | _0361_;
  assign _0522_ = ~_temp618_;
  assign _temp619_ = _0521_ & _0519_;
  assign _temp620_ = _temp619_ | _0522_;
  assign _0523_ = ~_temp620_;
  assign _0524_ = _0372_ & _0371_;
  assign _temp621_ = _0374_ & _0373_;
  assign _temp622_ = _temp621_ | _0524_;
  assign _0525_ = ~_temp622_;
  assign _0526_ = b[15] & a[7];
  assign _0527_ = b[16] & a[6];
  assign _0528_ = _0527_ ^ _0526_;
  assign _0529_ = b[17] & a[5];
  assign _temp623_ = _0529_ ^ _0528_;
  assign _0530_ = ~_temp623_;
  assign _0532_ = _0530_ ^ _0525_;
  assign _0533_ = _0396_ & _0395_;
  assign _0534_ = _0398_ & _0397_;
  assign _0535_ = _0534_ | _0533_;
  assign _temp624_ = _0535_ ^ _0532_;
  assign _0536_ = ~_temp624_;
  assign _temp625_ = _0399_ | _0394_;
  assign _0537_ = ~_temp625_;
  assign _temp626_ = _0404_ & _0400_;
  assign _temp627_ = _temp626_ | _0537_;
  assign _0538_ = ~_temp627_;
  assign _0539_ = _0538_ ^ _0536_;
  assign _0540_ = b[18] & a[4];
  assign _0541_ = b[19] & a[3];
  assign _0543_ = _0541_ ^ _0540_;
  assign _0544_ = b[20] & a[2];
  assign _temp628_ = _0544_ ^ _0543_;
  assign _0545_ = ~_temp628_;
  assign _0546_ = _0410_ & _0409_;
  assign _temp629_ = _0412_ & _0411_;
  assign _temp630_ = _temp629_ | _0546_;
  assign _0547_ = ~_temp630_;
  assign _temp631_ = _0547_ ^ _0545_;
  assign _0548_ = ~_temp631_;
  assign _temp632_ = b[21] & a[1];
  assign _0549_ = ~_temp632_;
  assign _0550_ = b[22] & a[0];
  assign _0551_ = _0550_ ^ _0549_;
  assign _0552_ = ~_0551_;
  assign _0554_ = _0552_ ^ _0548_;
  assign _0555_ = _0554_ ^ _0539_;
  assign _0556_ = _0555_ ^ _0523_;
  assign _temp633_ = _0407_ | _0405_;
  assign _0557_ = ~_temp633_;
  assign _0558_ = ~_0418_;
  assign _0559_ = _0558_ & _0408_;
  assign _0560_ = _0559_ | _0557_;
  assign _0561_ = _0560_ ^ _0556_;
  assign _temp634_ = _0561_ ^ _0518_;
  assign _0562_ = ~_temp634_;
  assign _temp635_ = _0386_ | _0384_;
  assign _0563_ = ~_temp635_;
  assign _temp636_ = _0426_ & _0387_;
  assign _temp637_ = _temp636_ | _0563_;
  assign _0565_ = ~_temp637_;
  assign _0566_ = _0565_ ^ _0562_;
  assign _temp638_ = _0419_ | _0392_;
  assign _0567_ = ~_temp638_;
  assign _0568_ = _0425_ & _0420_;
  assign _temp639_ = _0568_ | _0567_;
  assign _0569_ = ~_temp639_;
  assign _0570_ = ~_0416_;
  assign _temp640_ = _0415_ | _0413_;
  assign _0571_ = ~_temp640_;
  assign _temp641_ = _0417_ & _0570_;
  assign _temp642_ = _temp641_ | _0571_;
  assign _0572_ = ~_temp642_;
  assign _0573_ = _0572_ ^ _0569_;
  assign _temp643_ = _0573_ ^ _0566_;
  assign _0574_ = ~_temp643_;
  assign _temp644_ = _0429_ | _0427_;
  assign _0576_ = ~_temp644_;
  assign _temp645_ = _0438_ & _0430_;
  assign _temp646_ = _temp645_ | _0576_;
  assign _0577_ = ~_temp646_;
  assign _0578_ = _0577_ ^ _0574_;
  assign _0579_ = _0437_ & _0435_;
  assign _0580_ = _0579_ ^ _0578_;
  assign _temp647_ = _0441_ | _0439_;
  assign _0581_ = ~_temp647_;
  assign _0582_ = _0581_ ^ _0580_;
  assign _0583_ = _0443_ & _0442_;
  assign _0584_ = _0583_ ^ _0582_;
  assign _0585_ = _0446_ & _0445_;
  assign _temp648_ = _0448_ & _0447_;
  assign _temp649_ = _temp648_ | _0585_;
  assign _0587_ = ~_temp649_;
  assign _temp650_ = _0446_ ^ _0445_;
  assign _0588_ = ~_temp650_;
  assign _0589_ = _0588_ | _0310_;
  assign _temp651_ = _0589_ | _0319_;
  assign _temp652_ = _temp651_ & _0587_;
  assign _0590_ = ~_temp652_;
  assign q[22] = _0590_ ^ _0584_;
  assign _0591_ = a[23] & b[0];
  assign _0592_ = b[1] & a[22];
  assign _0593_ = _0592_ ^ _0591_;
  assign _0594_ = b[2] & a[21];
  assign _temp653_ = _0594_ ^ _0593_;
  assign _0595_ = ~_temp653_;
  assign _0597_ = _0452_ & _0451_;
  assign _temp654_ = _0455_ & _0453_;
  assign _temp655_ = _temp654_ | _0597_;
  assign _0598_ = ~_temp655_;
  assign _0599_ = _0598_ ^ _0595_;
  assign _0600_ = b[3] & a[20];
  assign _0601_ = b[4] & a[19];
  assign _0602_ = _0601_ ^ _0600_;
  assign _0603_ = b[5] & a[18];
  assign _0604_ = _0603_ ^ _0602_;
  assign _temp656_ = _0604_ ^ _0599_;
  assign _0605_ = ~_temp656_;
  assign _temp657_ = _0458_ | _0456_;
  assign _0606_ = ~_temp657_;
  assign _temp658_ = _0464_ & _0459_;
  assign _temp659_ = _temp658_ | _0606_;
  assign _0608_ = ~_temp659_;
  assign _0609_ = _0608_ ^ _0605_;
  assign _0610_ = _0461_ & _0460_;
  assign _0611_ = _0463_ & _0462_;
  assign _temp660_ = _0611_ | _0610_;
  assign _0612_ = ~_temp660_;
  assign _0613_ = b[6] & a[17];
  assign _0614_ = b[7] & a[16];
  assign _0615_ = _0614_ ^ _0613_;
  assign _0616_ = b[8] & a[15];
  assign _temp661_ = _0616_ ^ _0615_;
  assign _0617_ = ~_temp661_;
  assign _0619_ = _0617_ ^ _0612_;
  assign _0620_ = _0474_ & _0473_;
  assign _0621_ = _0477_ & _0475_;
  assign _0622_ = _0621_ | _0620_;
  assign _0623_ = _0622_ ^ _0619_;
  assign _temp662_ = _0623_ ^ _0609_;
  assign _0624_ = ~_temp662_;
  assign _temp663_ = _0468_ | _0466_;
  assign _0625_ = ~_temp663_;
  assign _temp664_ = _0483_ & _0469_;
  assign _temp665_ = _temp664_ | _0625_;
  assign _0626_ = ~_temp665_;
  assign _0627_ = _0626_ ^ _0624_;
  assign _temp666_ = _0478_ | _0472_;
  assign _0628_ = ~_temp666_;
  assign _temp667_ = _0482_ & _0479_;
  assign _temp668_ = _temp667_ | _0628_;
  assign _0630_ = ~_temp668_;
  assign _0631_ = b[9] & a[14];
  assign _0632_ = b[10] & a[13];
  assign _0633_ = _0632_ ^ _0631_;
  assign _0634_ = b[11] & a[12];
  assign _temp669_ = _0634_ ^ _0633_;
  assign _0635_ = ~_temp669_;
  assign _0636_ = _0494_ & _0493_;
  assign _temp670_ = _0496_ & _0495_;
  assign _temp671_ = _temp670_ | _0636_;
  assign _0637_ = ~_temp671_;
  assign _0638_ = _0637_ ^ _0635_;
  assign _0639_ = b[12] & a[11];
  assign _0641_ = b[13] & a[10];
  assign _0642_ = _0641_ ^ _0639_;
  assign _0643_ = b[14] & a[9];
  assign _temp672_ = _0643_ ^ _0642_;
  assign _0644_ = ~_temp672_;
  assign _0645_ = _0644_ ^ _0638_;
  assign _0646_ = _0645_ ^ _0630_;
  assign _temp673_ = _0500_ | _0497_;
  assign _0647_ = ~_temp673_;
  assign _0648_ = ~_0506_;
  assign _0649_ = _0648_ & _0501_;
  assign _0650_ = _0649_ | _0647_;
  assign _0652_ = _0650_ ^ _0646_;
  assign _temp674_ = _0652_ ^ _0627_;
  assign _0653_ = ~_temp674_;
  assign _temp675_ = _0486_ | _0484_;
  assign _0654_ = ~_temp675_;
  assign _temp676_ = _0514_ & _0488_;
  assign _temp677_ = _temp676_ | _0654_;
  assign _0655_ = ~_temp677_;
  assign _0656_ = _0655_ ^ _0653_;
  assign _temp678_ = _0507_ | _0492_;
  assign _0657_ = ~_temp678_;
  assign _temp679_ = _0513_ & _0508_;
  assign _temp680_ = _temp679_ | _0657_;
  assign _0658_ = ~_temp680_;
  assign _0659_ = _0503_ & _0502_;
  assign _0660_ = _0505_ & _0504_;
  assign _temp681_ = _0660_ | _0659_;
  assign _0661_ = ~_temp681_;
  assign _temp682_ = b[15] & a[8];
  assign _0663_ = ~_temp682_;
  assign _0664_ = b[16] & a[7];
  assign _0665_ = _0664_ ^ _0663_;
  assign _0666_ = b[17] & a[6];
  assign _0667_ = _0666_ ^ _0665_;
  assign _0668_ = _0667_ ^ _0661_;
  assign _0669_ = _0527_ & _0526_;
  assign _0670_ = _0529_ & _0528_;
  assign _0671_ = _0670_ | _0669_;
  assign _temp683_ = _0671_ ^ _0668_;
  assign _0672_ = ~_temp683_;
  assign _temp684_ = _0530_ | _0525_;
  assign _0673_ = ~_temp684_;
  assign _temp685_ = _0535_ & _0532_;
  assign _temp686_ = _temp685_ | _0673_;
  assign _0674_ = ~_temp686_;
  assign _0675_ = _0674_ ^ _0672_;
  assign _0676_ = b[18] & a[5];
  assign _0677_ = b[19] & a[4];
  assign _0678_ = _0677_ ^ _0676_;
  assign _0679_ = b[20] & a[3];
  assign _temp687_ = _0679_ ^ _0678_;
  assign _0680_ = ~_temp687_;
  assign _0681_ = _0541_ & _0540_;
  assign _temp688_ = _0544_ & _0543_;
  assign _temp689_ = _temp688_ | _0681_;
  assign _0682_ = ~_temp689_;
  assign _temp690_ = _0682_ ^ _0680_;
  assign _0684_ = ~_temp690_;
  assign _temp691_ = b[21] & a[2];
  assign _0685_ = ~_temp691_;
  assign _0686_ = b[22] & a[1];
  assign _0687_ = _0686_ ^ _0685_;
  assign _0688_ = b[23] & a[0];
  assign _0689_ = _0688_ ^ _0687_;
  assign _temp692_ = _0689_ ^ _0684_;
  assign _0690_ = ~_temp692_;
  assign _0691_ = _0690_ ^ _0675_;
  assign _0692_ = _0691_ ^ _0658_;
  assign _temp693_ = _0538_ | _0536_;
  assign _0693_ = ~_temp693_;
  assign _0695_ = ~_0554_;
  assign _0696_ = _0695_ & _0539_;
  assign _temp694_ = _0696_ | _0693_;
  assign _0697_ = ~_temp694_;
  assign _0698_ = ~_0697_;
  assign _0699_ = _0698_ ^ _0692_;
  assign _temp695_ = _0699_ ^ _0656_;
  assign _0700_ = ~_temp695_;
  assign _temp696_ = _0517_ | _0515_;
  assign _0701_ = ~_temp696_;
  assign _temp697_ = _0561_ & _0518_;
  assign _temp698_ = _temp697_ | _0701_;
  assign _0702_ = ~_temp698_;
  assign _0703_ = _0702_ ^ _0700_;
  assign _temp699_ = _0555_ | _0523_;
  assign _0704_ = ~_temp699_;
  assign _0706_ = _0560_ & _0556_;
  assign _temp700_ = _0706_ | _0704_;
  assign _0707_ = ~_temp700_;
  assign _temp701_ = _0547_ | _0545_;
  assign _0708_ = ~_temp701_;
  assign _temp702_ = _0551_ | _0548_;
  assign _0709_ = ~_temp702_;
  assign _temp703_ = _0709_ | _0708_;
  assign _0710_ = ~_temp703_;
  assign _0711_ = ~_0549_;
  assign _0712_ = _0550_ & _0711_;
  assign _0713_ = _0712_ ^ _0710_;
  assign _0714_ = _0713_ ^ _0707_;
  assign _temp704_ = _0714_ ^ _0703_;
  assign _0715_ = ~_temp704_;
  assign _temp705_ = _0565_ | _0562_;
  assign _0717_ = ~_temp705_;
  assign _temp706_ = _0573_ & _0566_;
  assign _temp707_ = _temp706_ | _0717_;
  assign _0718_ = ~_temp707_;
  assign _0719_ = _0718_ ^ _0715_;
  assign _temp708_ = _0572_ | _0569_;
  assign _0720_ = ~_temp708_;
  assign _temp709_ = _0720_ ^ _0719_;
  assign _0721_ = ~_temp709_;
  assign _temp710_ = _0577_ | _0574_;
  assign _0722_ = ~_temp710_;
  assign _temp711_ = _0579_ & _0578_;
  assign _temp712_ = _temp711_ | _0722_;
  assign _0723_ = ~_temp712_;
  assign _0724_ = _0723_ ^ _0721_;
  assign _0725_ = _0581_ & _0580_;
  assign _0726_ = _0725_ ^ _0724_;
  assign _0728_ = _0583_ & _0582_;
  assign _temp713_ = _0590_ & _0584_;
  assign _temp714_ = _temp713_ | _0728_;
  assign _0729_ = ~_temp714_;
  assign _temp715_ = _0729_ ^ _0726_;
  assign q[23] = ~_temp715_;
  assign _0730_ = a[24] & b[0];
  assign _0731_ = b[1] & a[23];
  assign _0732_ = _0731_ ^ _0730_;
  assign _0733_ = b[2] & a[22];
  assign _temp716_ = _0733_ ^ _0732_;
  assign _0734_ = ~_temp716_;
  assign _0735_ = _0592_ & _0591_;
  assign _temp717_ = _0594_ & _0593_;
  assign _temp718_ = _temp717_ | _0735_;
  assign _0736_ = ~_temp718_;
  assign _0738_ = _0736_ ^ _0734_;
  assign _0739_ = b[3] & a[21];
  assign _0740_ = b[4] & a[20];
  assign _0741_ = _0740_ ^ _0739_;
  assign _0742_ = b[5] & a[19];
  assign _temp719_ = _0742_ ^ _0741_;
  assign _0743_ = ~_temp719_;
  assign _0744_ = _0743_ ^ _0738_;
  assign _temp720_ = _0598_ | _0595_;
  assign _0745_ = ~_temp720_;
  assign _temp721_ = _0604_ & _0599_;
  assign _temp722_ = _temp721_ | _0745_;
  assign _0746_ = ~_temp722_;
  assign _0747_ = _0746_ ^ _0744_;
  assign _0749_ = _0601_ & _0600_;
  assign _0750_ = _0603_ & _0602_;
  assign _temp723_ = _0750_ | _0749_;
  assign _0751_ = ~_temp723_;
  assign _0752_ = b[6] & a[18];
  assign _0753_ = b[7] & a[17];
  assign _0754_ = _0753_ ^ _0752_;
  assign _0755_ = b[8] & a[16];
  assign _temp724_ = _0755_ ^ _0754_;
  assign _0756_ = ~_temp724_;
  assign _0757_ = _0756_ ^ _0751_;
  assign _0758_ = _0614_ & _0613_;
  assign _0760_ = _0616_ & _0615_;
  assign _0761_ = _0760_ | _0758_;
  assign _0762_ = _0761_ ^ _0757_;
  assign _temp725_ = _0762_ ^ _0747_;
  assign _0763_ = ~_temp725_;
  assign _temp726_ = _0608_ | _0605_;
  assign _0764_ = ~_temp726_;
  assign _temp727_ = _0623_ & _0609_;
  assign _temp728_ = _temp727_ | _0764_;
  assign _0765_ = ~_temp728_;
  assign _0766_ = _0765_ ^ _0763_;
  assign _temp729_ = _0617_ | _0612_;
  assign _0767_ = ~_temp729_;
  assign _0768_ = _0622_ & _0619_;
  assign _temp730_ = _0768_ | _0767_;
  assign _0769_ = ~_temp730_;
  assign _0771_ = b[9] & a[15];
  assign _0772_ = b[10] & a[14];
  assign _0773_ = _0772_ ^ _0771_;
  assign _0774_ = b[11] & a[13];
  assign _temp731_ = _0774_ ^ _0773_;
  assign _0775_ = ~_temp731_;
  assign _0776_ = _0632_ & _0631_;
  assign _temp732_ = _0634_ & _0633_;
  assign _temp733_ = _temp732_ | _0776_;
  assign _0777_ = ~_temp733_;
  assign _0778_ = _0777_ ^ _0775_;
  assign _0779_ = b[12] & a[12];
  assign _0780_ = b[13] & a[11];
  assign _0782_ = _0780_ ^ _0779_;
  assign _0783_ = b[14] & a[10];
  assign _temp734_ = _0783_ ^ _0782_;
  assign _0784_ = ~_temp734_;
  assign _0785_ = _0784_ ^ _0778_;
  assign _0786_ = _0785_ ^ _0769_;
  assign _temp735_ = _0637_ | _0635_;
  assign _0787_ = ~_temp735_;
  assign _0788_ = ~_0644_;
  assign _0789_ = _0788_ & _0638_;
  assign _temp736_ = _0789_ | _0787_;
  assign _0790_ = ~_temp736_;
  assign _0791_ = ~_0790_;
  assign _0793_ = _0791_ ^ _0786_;
  assign _temp737_ = _0793_ ^ _0766_;
  assign _0794_ = ~_temp737_;
  assign _temp738_ = _0626_ | _0624_;
  assign _0795_ = ~_temp738_;
  assign _temp739_ = _0652_ & _0627_;
  assign _temp740_ = _temp739_ | _0795_;
  assign _0796_ = ~_temp740_;
  assign _0797_ = _0796_ ^ _0794_;
  assign _temp741_ = _0645_ | _0630_;
  assign _0798_ = ~_temp741_;
  assign _0799_ = _0650_ & _0646_;
  assign _temp742_ = _0799_ | _0798_;
  assign _0800_ = ~_temp742_;
  assign _0801_ = _0641_ & _0639_;
  assign _temp743_ = _0643_ & _0642_;
  assign _temp744_ = _temp743_ | _0801_;
  assign _0802_ = ~_temp744_;
  assign _0804_ = b[15] & a[9];
  assign _0805_ = b[16] & a[8];
  assign _temp745_ = _0805_ ^ _0804_;
  assign _0806_ = ~_temp745_;
  assign _0807_ = b[17] & a[7];
  assign _0808_ = _0807_ ^ _0806_;
  assign _0809_ = _0808_ ^ _0802_;
  assign _0810_ = ~_0663_;
  assign _0811_ = _0664_ & _0810_;
  assign _0812_ = ~_0666_;
  assign _temp746_ = _0812_ | _0665_;
  assign _0813_ = ~_temp746_;
  assign _temp747_ = _0813_ | _0811_;
  assign _0815_ = ~_temp747_;
  assign _0816_ = _0815_ ^ _0809_;
  assign _temp748_ = _0667_ | _0661_;
  assign _0817_ = ~_temp748_;
  assign _temp749_ = _0671_ & _0668_;
  assign _temp750_ = _temp749_ | _0817_;
  assign _0818_ = ~_temp750_;
  assign _0819_ = _0818_ ^ _0816_;
  assign _0820_ = b[18] & a[6];
  assign _0821_ = b[19] & a[5];
  assign _0822_ = _0821_ ^ _0820_;
  assign _0823_ = b[20] & a[4];
  assign _temp751_ = _0823_ ^ _0822_;
  assign _0824_ = ~_temp751_;
  assign _0826_ = _0677_ & _0676_;
  assign _temp752_ = _0679_ & _0678_;
  assign _temp753_ = _temp752_ | _0826_;
  assign _0827_ = ~_temp753_;
  assign _temp754_ = _0827_ ^ _0824_;
  assign _0828_ = ~_temp754_;
  assign _0829_ = b[21] & a[3];
  assign _0830_ = b[22] & a[2];
  assign _temp755_ = _0830_ ^ _0829_;
  assign _0831_ = ~_temp755_;
  assign _0832_ = b[23] & a[1];
  assign _0833_ = _0832_ ^ _0831_;
  assign _0834_ = ~_0833_;
  assign _0835_ = _0834_ ^ _0828_;
  assign _0837_ = _0835_ ^ _0819_;
  assign _0838_ = _0837_ ^ _0800_;
  assign _temp756_ = _0674_ | _0672_;
  assign _0839_ = ~_temp756_;
  assign _0840_ = ~_0690_;
  assign _0841_ = _0840_ & _0675_;
  assign _0842_ = _0841_ | _0839_;
  assign _0843_ = _0842_ ^ _0838_;
  assign _temp757_ = _0843_ ^ _0797_;
  assign _0844_ = ~_temp757_;
  assign _temp758_ = _0655_ | _0653_;
  assign _0845_ = ~_temp758_;
  assign _temp759_ = _0699_ & _0656_;
  assign _temp760_ = _temp759_ | _0845_;
  assign _0846_ = ~_temp760_;
  assign _0848_ = _0846_ ^ _0844_;
  assign _temp761_ = _0691_ | _0658_;
  assign _0849_ = ~_temp761_;
  assign _0850_ = _0698_ & _0692_;
  assign _temp762_ = _0850_ | _0849_;
  assign _0851_ = ~_temp762_;
  assign _0852_ = _0682_ | _0680_;
  assign _temp763_ = _0689_ | _0684_;
  assign _temp764_ = _temp763_ & _0852_;
  assign _0853_ = ~_temp764_;
  assign _0854_ = ~_0685_;
  assign _0855_ = _0686_ & _0854_;
  assign _0856_ = ~_0688_;
  assign _temp765_ = _0856_ | _0687_;
  assign _0857_ = ~_temp765_;
  assign _temp766_ = _0857_ | _0855_;
  assign _0859_ = ~_temp766_;
  assign _0860_ = a[0] & b[24];
  assign _0861_ = _0860_ ^ _0859_;
  assign _0862_ = _0861_ ^ _0853_;
  assign _0863_ = ~_0712_;
  assign _temp767_ = _0863_ | _0710_;
  assign _0864_ = ~_temp767_;
  assign _0865_ = _0864_ ^ _0862_;
  assign _0866_ = _0865_ ^ _0851_;
  assign _temp768_ = _0866_ ^ _0848_;
  assign _0867_ = ~_temp768_;
  assign _temp769_ = _0702_ | _0700_;
  assign _0868_ = ~_temp769_;
  assign _temp770_ = _0714_ & _0703_;
  assign _temp771_ = _temp770_ | _0868_;
  assign _0870_ = ~_temp771_;
  assign _0871_ = _0870_ ^ _0867_;
  assign _temp772_ = _0713_ | _0707_;
  assign _0872_ = ~_temp772_;
  assign _temp773_ = _0872_ ^ _0871_;
  assign _0873_ = ~_temp773_;
  assign _temp774_ = _0718_ | _0715_;
  assign _0874_ = ~_temp774_;
  assign _temp775_ = _0720_ & _0719_;
  assign _temp776_ = _temp775_ | _0874_;
  assign _0875_ = ~_temp776_;
  assign _0876_ = _0875_ ^ _0873_;
  assign _temp777_ = _0723_ | _0721_;
  assign _0877_ = ~_temp777_;
  assign _0878_ = _0877_ ^ _0876_;
  assign _temp778_ = _0726_ & _0584_;
  assign _0879_ = ~_temp778_;
  assign _0881_ = _0879_ | _0589_;
  assign _temp779_ = _0879_ | _0589_;
  assign _0882_ = ~_temp779_;
  assign _0883_ = _0725_ & _0724_;
  assign _temp780_ = _0728_ & _0726_;
  assign _temp781_ = _temp780_ | _0883_;
  assign _0884_ = ~_temp781_;
  assign _temp782_ = _0879_ | _0587_;
  assign _temp783_ = _temp782_ & _0884_;
  assign _0885_ = ~_temp783_;
  assign _temp784_ = _0882_ & _0315_;
  assign _temp785_ = _temp784_ | _0885_;
  assign _0886_ = ~_temp785_;
  assign _temp786_ = _0881_ | _0318_;
  assign _temp787_ = _temp786_ & _0886_;
  assign _0887_ = ~_temp787_;
  assign q[24] = _0887_ ^ _0878_;
  assign _0888_ = a[25] & b[0];
  assign _0889_ = b[1] & a[24];
  assign _0891_ = _0889_ ^ _0888_;
  assign _0892_ = b[2] & a[23];
  assign _temp788_ = _0892_ ^ _0891_;
  assign _0893_ = ~_temp788_;
  assign _0894_ = _0731_ & _0730_;
  assign _temp789_ = _0733_ & _0732_;
  assign _temp790_ = _temp789_ | _0894_;
  assign _0895_ = ~_temp790_;
  assign _0896_ = _0895_ ^ _0893_;
  assign _0897_ = b[3] & a[22];
  assign _0898_ = b[4] & a[21];
  assign _0899_ = _0898_ ^ _0897_;
  assign _0900_ = b[5] & a[20];
  assign _temp791_ = _0900_ ^ _0899_;
  assign _0902_ = ~_temp791_;
  assign _0903_ = _0902_ ^ _0896_;
  assign _0904_ = ~_0743_;
  assign _temp792_ = _0736_ | _0734_;
  assign _0905_ = ~_temp792_;
  assign _temp793_ = _0904_ & _0738_;
  assign _temp794_ = _temp793_ | _0905_;
  assign _0906_ = ~_temp794_;
  assign _temp795_ = _0906_ ^ _0903_;
  assign _0907_ = ~_temp795_;
  assign _0908_ = _0740_ & _0739_;
  assign _0909_ = _0742_ & _0741_;
  assign _temp796_ = _0909_ | _0908_;
  assign _0910_ = ~_temp796_;
  assign _temp797_ = b[6] & a[19];
  assign _0911_ = ~_temp797_;
  assign _0913_ = b[7] & a[18];
  assign _0914_ = _0913_ ^ _0911_;
  assign _0915_ = b[8] & a[17];
  assign _0916_ = _0915_ ^ _0914_;
  assign _0917_ = _0916_ ^ _0910_;
  assign _0918_ = _0753_ & _0752_;
  assign _0919_ = _0755_ & _0754_;
  assign _0920_ = _0919_ | _0918_;
  assign _temp798_ = _0920_ ^ _0917_;
  assign _0921_ = ~_temp798_;
  assign _temp799_ = _0921_ ^ _0907_;
  assign _0922_ = ~_temp799_;
  assign _temp800_ = _0746_ | _0744_;
  assign _0924_ = ~_temp800_;
  assign _temp801_ = _0762_ & _0747_;
  assign _temp802_ = _temp801_ | _0924_;
  assign _0925_ = ~_temp802_;
  assign _temp803_ = _0925_ ^ _0922_;
  assign _0926_ = ~_temp803_;
  assign _0927_ = ~_0926_;
  assign _temp804_ = _0756_ | _0751_;
  assign _0928_ = ~_temp804_;
  assign _0929_ = _0761_ & _0757_;
  assign _temp805_ = _0929_ | _0928_;
  assign _0930_ = ~_temp805_;
  assign _0931_ = b[9] & a[16];
  assign _0932_ = b[10] & a[15];
  assign _0933_ = _0932_ ^ _0931_;
  assign _0935_ = b[11] & a[14];
  assign _temp806_ = _0935_ ^ _0933_;
  assign _0936_ = ~_temp806_;
  assign _0937_ = _0772_ & _0771_;
  assign _temp807_ = _0774_ & _0773_;
  assign _temp808_ = _temp807_ | _0937_;
  assign _0938_ = ~_temp808_;
  assign _0939_ = _0938_ ^ _0936_;
  assign _0940_ = b[12] & a[13];
  assign _0941_ = b[13] & a[12];
  assign _0942_ = _0941_ ^ _0940_;
  assign _0943_ = b[14] & a[11];
  assign _temp809_ = _0943_ ^ _0942_;
  assign _0944_ = ~_temp809_;
  assign _0946_ = _0944_ ^ _0939_;
  assign _0947_ = _0946_ ^ _0930_;
  assign _temp810_ = _0777_ | _0775_;
  assign _0948_ = ~_temp810_;
  assign _0949_ = ~_0784_;
  assign _0950_ = _0949_ & _0778_;
  assign _temp811_ = _0950_ | _0948_;
  assign _0951_ = ~_temp811_;
  assign _0952_ = _0951_ ^ _0947_;
  assign _0953_ = _0952_ ^ _0927_;
  assign _temp812_ = _0765_ | _0763_;
  assign _0954_ = ~_temp812_;
  assign _temp813_ = _0793_ & _0766_;
  assign _temp814_ = _temp813_ | _0954_;
  assign _0955_ = ~_temp814_;
  assign _0957_ = _0955_ ^ _0953_;
  assign _temp815_ = _0785_ | _0769_;
  assign _0958_ = ~_temp815_;
  assign _0959_ = _0791_ & _0786_;
  assign _temp816_ = _0959_ | _0958_;
  assign _0960_ = ~_temp816_;
  assign _0961_ = _0780_ & _0779_;
  assign _temp817_ = _0783_ & _0782_;
  assign _temp818_ = _temp817_ | _0961_;
  assign _0962_ = ~_temp818_;
  assign _0963_ = b[15] & a[10];
  assign _0964_ = b[16] & a[9];
  assign _temp819_ = _0964_ ^ _0963_;
  assign _0965_ = ~_temp819_;
  assign _0966_ = b[17] & a[8];
  assign _0968_ = _0966_ ^ _0965_;
  assign _0969_ = _0968_ ^ _0962_;
  assign _0970_ = _0805_ & _0804_;
  assign _0971_ = ~_0807_;
  assign _temp820_ = _0971_ | _0806_;
  assign _0972_ = ~_temp820_;
  assign _temp821_ = _0972_ | _0970_;
  assign _0973_ = ~_temp821_;
  assign _0974_ = _0973_ ^ _0969_;
  assign _0975_ = ~_0815_;
  assign _temp822_ = _0808_ | _0802_;
  assign _0976_ = ~_temp822_;
  assign _temp823_ = _0975_ & _0809_;
  assign _temp824_ = _temp823_ | _0976_;
  assign _0977_ = ~_temp824_;
  assign _0979_ = _0977_ ^ _0974_;
  assign _0980_ = b[18] & a[7];
  assign _0981_ = b[19] & a[6];
  assign _0982_ = _0981_ ^ _0980_;
  assign _0983_ = b[20] & a[5];
  assign _temp825_ = _0983_ ^ _0982_;
  assign _0984_ = ~_temp825_;
  assign _0985_ = _0821_ & _0820_;
  assign _temp826_ = _0823_ & _0822_;
  assign _temp827_ = _temp826_ | _0985_;
  assign _0986_ = ~_temp827_;
  assign _0987_ = _0986_ ^ _0984_;
  assign _0988_ = b[21] & a[4];
  assign _0990_ = b[22] & a[3];
  assign _0991_ = _0990_ ^ _0988_;
  assign _0992_ = b[23] & a[2];
  assign _temp828_ = _0992_ ^ _0991_;
  assign _0993_ = ~_temp828_;
  assign _0994_ = _0993_ ^ _0987_;
  assign _0995_ = _0994_ ^ _0979_;
  assign _temp829_ = _0995_ ^ _0960_;
  assign _0996_ = ~_temp829_;
  assign _temp830_ = _0818_ | _0816_;
  assign _0997_ = ~_temp830_;
  assign _0998_ = ~_0835_;
  assign _0999_ = _0998_ & _0819_;
  assign _temp831_ = _0999_ | _0997_;
  assign _1001_ = ~_temp831_;
  assign _1002_ = _1001_ ^ _0996_;
  assign _temp832_ = _1002_ ^ _0957_;
  assign _1003_ = ~_temp832_;
  assign _temp833_ = _0796_ | _0794_;
  assign _1004_ = ~_temp833_;
  assign _temp834_ = _0843_ & _0797_;
  assign _temp835_ = _temp834_ | _1004_;
  assign _1005_ = ~_temp835_;
  assign _1006_ = _1005_ ^ _1003_;
  assign _temp836_ = _0837_ | _0800_;
  assign _1007_ = ~_temp836_;
  assign _1008_ = _0842_ & _0838_;
  assign _temp837_ = _1008_ | _1007_;
  assign _1009_ = ~_temp837_;
  assign _temp838_ = _0827_ | _0824_;
  assign _1010_ = ~_temp838_;
  assign _temp839_ = _0833_ | _0828_;
  assign _1012_ = ~_temp839_;
  assign _temp840_ = _1012_ | _1010_;
  assign _1013_ = ~_temp840_;
  assign _1014_ = _0830_ & _0829_;
  assign _1015_ = ~_0832_;
  assign _temp841_ = _1015_ | _0831_;
  assign _1016_ = ~_temp841_;
  assign _temp842_ = _1016_ | _1014_;
  assign _1017_ = ~_temp842_;
  assign _1018_ = a[1] & b[24];
  assign _1019_ = b[25] & a[0];
  assign _temp843_ = _1019_ ^ _1018_;
  assign _1020_ = ~_temp843_;
  assign _temp844_ = _1020_ ^ _1017_;
  assign _1021_ = ~_temp844_;
  assign _temp845_ = _1021_ ^ _1013_;
  assign _1022_ = ~_temp845_;
  assign _1023_ = ~_0860_;
  assign _temp846_ = _1023_ | _0859_;
  assign _1024_ = ~_temp846_;
  assign _1025_ = _1024_ ^ _1022_;
  assign _1026_ = ~_0861_;
  assign _1027_ = _1026_ & _0853_;
  assign _1028_ = _1027_ ^ _1025_;
  assign _1029_ = _1028_ ^ _1009_;
  assign _1030_ = ~_0862_;
  assign _1031_ = _0864_ & _1030_;
  assign _1033_ = _1031_ ^ _1029_;
  assign _temp847_ = _1033_ ^ _1006_;
  assign _1034_ = ~_temp847_;
  assign _temp848_ = _0846_ | _0844_;
  assign _1035_ = ~_temp848_;
  assign _temp849_ = _0866_ & _0848_;
  assign _temp850_ = _temp849_ | _1035_;
  assign _1036_ = ~_temp850_;
  assign _1037_ = _1036_ ^ _1034_;
  assign _temp851_ = _0865_ | _0851_;
  assign _1038_ = ~_temp851_;
  assign _temp852_ = _1038_ ^ _1037_;
  assign _1039_ = ~_temp852_;
  assign _temp853_ = _0870_ | _0867_;
  assign _1040_ = ~_temp853_;
  assign _temp854_ = _0872_ & _0871_;
  assign _temp855_ = _temp854_ | _1040_;
  assign _1041_ = ~_temp855_;
  assign _1042_ = _1041_ ^ _1039_;
  assign _temp856_ = _0875_ | _0873_;
  assign _1044_ = ~_temp856_;
  assign _1045_ = _1044_ ^ _1042_;
  assign _1046_ = _0877_ & _0876_;
  assign _temp857_ = _0887_ & _0878_;
  assign _temp858_ = _temp857_ | _1046_;
  assign _1047_ = ~_temp858_;
  assign _temp859_ = _1047_ ^ _1045_;
  assign q[25] = ~_temp859_;
  assign _1048_ = a[26] & b[0];
  assign _1049_ = b[1] & a[25];
  assign _1050_ = _1049_ ^ _1048_;
  assign _1051_ = b[2] & a[24];
  assign _temp860_ = _1051_ ^ _1050_;
  assign _1052_ = ~_temp860_;
  assign _1054_ = _0889_ & _0888_;
  assign _temp861_ = _0892_ & _0891_;
  assign _temp862_ = _temp861_ | _1054_;
  assign _1055_ = ~_temp862_;
  assign _1056_ = _1055_ ^ _1052_;
  assign _1057_ = b[3] & a[23];
  assign _1058_ = b[4] & a[22];
  assign _temp863_ = _1058_ ^ _1057_;
  assign _1059_ = ~_temp863_;
  assign _1060_ = b[5] & a[21];
  assign _1061_ = _1060_ ^ _1059_;
  assign _1062_ = _1061_ ^ _1056_;
  assign _1063_ = ~_0902_;
  assign _temp864_ = _0895_ | _0893_;
  assign _1065_ = ~_temp864_;
  assign _temp865_ = _1063_ & _0896_;
  assign _temp866_ = _temp865_ | _1065_;
  assign _1066_ = ~_temp866_;
  assign _1067_ = _1066_ ^ _1062_;
  assign _1068_ = _0898_ & _0897_;
  assign _1069_ = _0900_ & _0899_;
  assign _temp867_ = _1069_ | _1068_;
  assign _1070_ = ~_temp867_;
  assign _1071_ = b[6] & a[20];
  assign _1072_ = b[7] & a[19];
  assign _temp868_ = _1072_ ^ _1071_;
  assign _1073_ = ~_temp868_;
  assign _1074_ = b[8] & a[18];
  assign _1076_ = _1074_ ^ _1073_;
  assign _1077_ = _1076_ ^ _1070_;
  assign _1078_ = ~_0911_;
  assign _1079_ = _0913_ & _1078_;
  assign _1080_ = ~_0915_;
  assign _temp869_ = _1080_ | _0914_;
  assign _1081_ = ~_temp869_;
  assign _temp870_ = _1081_ | _1079_;
  assign _1082_ = ~_temp870_;
  assign _1083_ = _1082_ ^ _1077_;
  assign _1084_ = _1083_ ^ _1067_;
  assign _1085_ = _0906_ | _0903_;
  assign _1087_ = _0921_ | _0907_;
  assign _1088_ = _1087_ & _1085_;
  assign _1089_ = _1088_ ^ _1084_;
  assign _temp871_ = _0916_ | _0910_;
  assign _1090_ = ~_temp871_;
  assign _1091_ = _0920_ & _0917_;
  assign _temp872_ = _1091_ | _1090_;
  assign _1092_ = ~_temp872_;
  assign _1093_ = b[9] & a[17];
  assign _1094_ = b[10] & a[16];
  assign _temp873_ = _1094_ ^ _1093_;
  assign _1095_ = ~_temp873_;
  assign _1096_ = b[11] & a[15];
  assign _1098_ = _1096_ ^ _1095_;
  assign _1099_ = _0932_ & _0931_;
  assign _temp874_ = _0935_ & _0933_;
  assign _temp875_ = _temp874_ | _1099_;
  assign _1100_ = ~_temp875_;
  assign _1101_ = _1100_ ^ _1098_;
  assign _1102_ = b[12] & a[14];
  assign _1103_ = b[13] & a[13];
  assign _temp876_ = _1103_ ^ _1102_;
  assign _1104_ = ~_temp876_;
  assign _1105_ = b[14] & a[12];
  assign _1106_ = _1105_ ^ _1104_;
  assign _1107_ = _1106_ ^ _1101_;
  assign _1109_ = _1107_ ^ _1092_;
  assign _temp877_ = _0938_ | _0936_;
  assign _1110_ = ~_temp877_;
  assign _1111_ = ~_0944_;
  assign _1112_ = _1111_ & _0939_;
  assign _temp878_ = _1112_ | _1110_;
  assign _1113_ = ~_temp878_;
  assign _1114_ = ~_1113_;
  assign _1115_ = _1114_ ^ _1109_;
  assign _temp879_ = _1115_ ^ _1089_;
  assign _1116_ = ~_temp879_;
  assign _1117_ = _0925_ | _0922_;
  assign _1118_ = _0952_ | _0926_;
  assign _1120_ = _1118_ & _1117_;
  assign _1121_ = _1120_ ^ _1116_;
  assign _temp880_ = _0946_ | _0930_;
  assign _1122_ = ~_temp880_;
  assign _1123_ = ~_0951_;
  assign _1124_ = _1123_ & _0947_;
  assign _temp881_ = _1124_ | _1122_;
  assign _1125_ = ~_temp881_;
  assign _1126_ = _0941_ & _0940_;
  assign _temp882_ = _0943_ & _0942_;
  assign _temp883_ = _temp882_ | _1126_;
  assign _1127_ = ~_temp883_;
  assign _1128_ = b[15] & a[11];
  assign _1129_ = b[16] & a[10];
  assign _temp884_ = _1129_ ^ _1128_;
  assign _1131_ = ~_temp884_;
  assign _1132_ = b[17] & a[9];
  assign _1133_ = _1132_ ^ _1131_;
  assign _1134_ = _1133_ ^ _1127_;
  assign _1135_ = _0964_ & _0963_;
  assign _1136_ = ~_0966_;
  assign _temp885_ = _1136_ | _0965_;
  assign _1137_ = ~_temp885_;
  assign _temp886_ = _1137_ | _1135_;
  assign _1138_ = ~_temp886_;
  assign _1139_ = _1138_ ^ _1134_;
  assign _1140_ = ~_0973_;
  assign _temp887_ = _0968_ | _0962_;
  assign _1142_ = ~_temp887_;
  assign _temp888_ = _1140_ & _0969_;
  assign _temp889_ = _temp888_ | _1142_;
  assign _1143_ = ~_temp889_;
  assign _1144_ = _1143_ ^ _1139_;
  assign _1145_ = b[18] & a[8];
  assign _1146_ = b[19] & a[7];
  assign _temp890_ = _1146_ ^ _1145_;
  assign _1147_ = ~_temp890_;
  assign _1148_ = b[20] & a[6];
  assign _1149_ = _1148_ ^ _1147_;
  assign _1150_ = _0981_ & _0980_;
  assign _temp891_ = _0983_ & _0982_;
  assign _temp892_ = _temp891_ | _1150_;
  assign _1151_ = ~_temp892_;
  assign _temp893_ = _1151_ ^ _1149_;
  assign _1153_ = ~_temp893_;
  assign _1154_ = b[21] & a[5];
  assign _1155_ = b[22] & a[4];
  assign _temp894_ = _1155_ ^ _1154_;
  assign _1156_ = ~_temp894_;
  assign _1157_ = b[23] & a[3];
  assign _1158_ = _1157_ ^ _1156_;
  assign _1159_ = ~_1158_;
  assign _1160_ = _1159_ ^ _1153_;
  assign _1161_ = _1160_ ^ _1144_;
  assign _temp895_ = _1161_ ^ _1125_;
  assign _1162_ = ~_temp895_;
  assign _1164_ = ~_0994_;
  assign _temp896_ = _0977_ | _0974_;
  assign _1165_ = ~_temp896_;
  assign _temp897_ = _1164_ & _0979_;
  assign _temp898_ = _temp897_ | _1165_;
  assign _1166_ = ~_temp898_;
  assign _1167_ = _1166_ ^ _1162_;
  assign _temp899_ = _1167_ ^ _1121_;
  assign _1168_ = ~_temp899_;
  assign _temp900_ = _0955_ | _0953_;
  assign _1169_ = ~_temp900_;
  assign _temp901_ = _1002_ & _0957_;
  assign _temp902_ = _temp901_ | _1169_;
  assign _1170_ = ~_temp902_;
  assign _1171_ = _1170_ ^ _1168_;
  assign _1172_ = _0995_ ^ _0960_;
  assign _1173_ = ~_1001_;
  assign _temp903_ = _0995_ | _0960_;
  assign _1175_ = ~_temp903_;
  assign _temp904_ = _1173_ & _1172_;
  assign _temp905_ = _temp904_ | _1175_;
  assign _1176_ = ~_temp905_;
  assign _temp906_ = _0986_ | _0984_;
  assign _1177_ = ~_temp906_;
  assign _1178_ = ~_0993_;
  assign _1179_ = _1178_ & _0987_;
  assign _temp907_ = _1179_ | _1177_;
  assign _1180_ = ~_temp907_;
  assign _1181_ = _0990_ & _0988_;
  assign _1182_ = _0992_ & _0991_;
  assign _1183_ = _1182_ | _1181_;
  assign _1184_ = a[2] & b[24];
  assign _1186_ = a[1] & b[25];
  assign _temp908_ = _1186_ ^ _1184_;
  assign _1187_ = ~_temp908_;
  assign _1188_ = b[26] & a[0];
  assign _1189_ = _1188_ ^ _1187_;
  assign _1190_ = _1189_ ^ _1183_;
  assign _1191_ = _1019_ & _1018_;
  assign _1192_ = _1191_ ^ _1190_;
  assign _1193_ = _1192_ ^ _1180_;
  assign _temp909_ = _1020_ | _1017_;
  assign _1194_ = ~_temp909_;
  assign _temp910_ = _1194_ ^ _1193_;
  assign _1195_ = ~_temp910_;
  assign _1197_ = ~_1022_;
  assign _temp911_ = _1021_ | _1013_;
  assign _1198_ = ~_temp911_;
  assign _temp912_ = _1024_ & _1197_;
  assign _temp913_ = _temp912_ | _1198_;
  assign _1199_ = ~_temp913_;
  assign _temp914_ = _1199_ ^ _1195_;
  assign _1200_ = ~_temp914_;
  assign _1201_ = _1200_ ^ _1176_;
  assign _1202_ = ~_1027_;
  assign _temp915_ = _1202_ | _1025_;
  assign _1203_ = ~_temp915_;
  assign _1204_ = _1203_ ^ _1201_;
  assign _temp916_ = _1204_ ^ _1171_;
  assign _1205_ = ~_temp916_;
  assign _temp917_ = _1005_ | _1003_;
  assign _1206_ = ~_temp917_;
  assign _temp918_ = _1033_ & _1006_;
  assign _temp919_ = _temp918_ | _1206_;
  assign _1208_ = ~_temp919_;
  assign _1209_ = _1208_ ^ _1205_;
  assign _temp920_ = _1028_ | _1009_;
  assign _1210_ = ~_temp920_;
  assign _1211_ = _1031_ & _1029_;
  assign _1212_ = _1211_ | _1210_;
  assign _temp921_ = _1212_ ^ _1209_;
  assign _1213_ = ~_temp921_;
  assign _temp922_ = _1036_ | _1034_;
  assign _1214_ = ~_temp922_;
  assign _temp923_ = _1038_ & _1037_;
  assign _temp924_ = _temp923_ | _1214_;
  assign _1215_ = ~_temp924_;
  assign _1216_ = _1215_ ^ _1213_;
  assign _temp925_ = _1041_ | _1039_;
  assign _1217_ = ~_temp925_;
  assign _1219_ = _1217_ ^ _1216_;
  assign _1220_ = _0881_ | _0318_;
  assign _1221_ = _0886_ & _1220_;
  assign _1222_ = _1044_ & _1042_;
  assign _temp926_ = _1046_ & _1045_;
  assign _temp927_ = _temp926_ | _1222_;
  assign _1223_ = ~_temp927_;
  assign _temp928_ = _1045_ & _0878_;
  assign _1224_ = ~_temp928_;
  assign _temp929_ = _1224_ | _1221_;
  assign _temp930_ = _temp929_ & _1223_;
  assign _1225_ = ~_temp930_;
  assign q[26] = _1225_ ^ _1219_;
  assign _1226_ = a[27] & b[0];
  assign _1227_ = b[1] & a[26];
  assign _temp931_ = _1227_ ^ _1226_;
  assign _1229_ = ~_temp931_;
  assign _1230_ = b[2] & a[25];
  assign _1231_ = _1230_ ^ _1229_;
  assign _1232_ = _1049_ & _1048_;
  assign _temp932_ = _1051_ & _1050_;
  assign _temp933_ = _temp932_ | _1232_;
  assign _1233_ = ~_temp933_;
  assign _temp934_ = _1233_ ^ _1231_;
  assign _1234_ = ~_temp934_;
  assign _temp935_ = b[3] & a[24];
  assign _1235_ = ~_temp935_;
  assign _1236_ = b[4] & a[23];
  assign _1237_ = _1236_ ^ _1235_;
  assign _1238_ = b[5] & a[22];
  assign _1240_ = _1238_ ^ _1237_;
  assign _1241_ = ~_1240_;
  assign _1242_ = _1241_ ^ _1234_;
  assign _1243_ = ~_1061_;
  assign _temp936_ = _1055_ | _1052_;
  assign _1244_ = ~_temp936_;
  assign _temp937_ = _1243_ & _1056_;
  assign _temp938_ = _temp937_ | _1244_;
  assign _1245_ = ~_temp938_;
  assign _temp939_ = _1245_ ^ _1242_;
  assign _1246_ = ~_temp939_;
  assign _1247_ = _1058_ & _1057_;
  assign _1248_ = ~_1060_;
  assign _temp940_ = _1248_ | _1059_;
  assign _1249_ = ~_temp940_;
  assign _temp941_ = _1249_ | _1247_;
  assign _1251_ = ~_temp941_;
  assign _temp942_ = b[6] & a[21];
  assign _1252_ = ~_temp942_;
  assign _1253_ = b[7] & a[20];
  assign _1254_ = _1253_ ^ _1252_;
  assign _1255_ = b[8] & a[19];
  assign _1256_ = _1255_ ^ _1254_;
  assign _temp943_ = _1256_ ^ _1251_;
  assign _1257_ = ~_temp943_;
  assign _1258_ = _1072_ & _1071_;
  assign _1259_ = ~_1074_;
  assign _temp944_ = _1259_ | _1073_;
  assign _1260_ = ~_temp944_;
  assign _temp945_ = _1260_ | _1258_;
  assign _1262_ = ~_temp945_;
  assign _1263_ = ~_1262_;
  assign _1264_ = _1263_ ^ _1257_;
  assign _temp946_ = _1264_ ^ _1246_;
  assign _1265_ = ~_temp946_;
  assign _1266_ = ~_1083_;
  assign _temp947_ = _1066_ | _1062_;
  assign _1267_ = ~_temp947_;
  assign _temp948_ = _1266_ & _1067_;
  assign _temp949_ = _temp948_ | _1267_;
  assign _1268_ = ~_temp949_;
  assign _1269_ = _1268_ ^ _1265_;
  assign _temp950_ = _1076_ | _1070_;
  assign _1270_ = ~_temp950_;
  assign _1271_ = ~_1082_;
  assign _1273_ = _1271_ & _1077_;
  assign _temp951_ = _1273_ | _1270_;
  assign _1274_ = ~_temp951_;
  assign _temp952_ = b[9] & a[18];
  assign _1275_ = ~_temp952_;
  assign _1276_ = b[10] & a[17];
  assign _1277_ = _1276_ ^ _1275_;
  assign _1278_ = b[11] & a[16];
  assign _1279_ = _1278_ ^ _1277_;
  assign _1280_ = ~_1095_;
  assign _1281_ = _1094_ & _1093_;
  assign _temp953_ = _1096_ & _1280_;
  assign _temp954_ = _temp953_ | _1281_;
  assign _1282_ = ~_temp954_;
  assign _1284_ = _1282_ ^ _1279_;
  assign _temp955_ = b[12] & a[15];
  assign _1285_ = ~_temp955_;
  assign _1286_ = b[13] & a[14];
  assign _1287_ = _1286_ ^ _1285_;
  assign _1288_ = b[14] & a[13];
  assign _1289_ = _1288_ ^ _1287_;
  assign _1290_ = _1289_ ^ _1284_;
  assign _1291_ = _1290_ ^ _1274_;
  assign _temp956_ = _1100_ | _1098_;
  assign _1292_ = ~_temp956_;
  assign _1293_ = ~_1106_;
  assign _1295_ = _1293_ & _1101_;
  assign _temp957_ = _1295_ | _1292_;
  assign _1296_ = ~_temp957_;
  assign _1297_ = ~_1296_;
  assign _1298_ = _1297_ ^ _1291_;
  assign _temp958_ = _1298_ ^ _1269_;
  assign _1299_ = ~_temp958_;
  assign _temp959_ = _1088_ | _1084_;
  assign _1300_ = ~_temp959_;
  assign _temp960_ = _1115_ & _1089_;
  assign _temp961_ = _temp960_ | _1300_;
  assign _1301_ = ~_temp961_;
  assign _1302_ = _1301_ ^ _1299_;
  assign _temp962_ = _1107_ | _1092_;
  assign _1303_ = ~_temp962_;
  assign _1304_ = _1114_ & _1109_;
  assign _temp963_ = _1304_ | _1303_;
  assign _1306_ = ~_temp963_;
  assign _1307_ = ~_1104_;
  assign _1308_ = _1103_ & _1102_;
  assign _temp964_ = _1105_ & _1307_;
  assign _temp965_ = _temp964_ | _1308_;
  assign _1309_ = ~_temp965_;
  assign _temp966_ = b[15] & a[12];
  assign _1310_ = ~_temp966_;
  assign _1311_ = b[16] & a[11];
  assign _1312_ = _1311_ ^ _1310_;
  assign _1313_ = b[17] & a[10];
  assign _1314_ = _1313_ ^ _1312_;
  assign _1315_ = _1314_ ^ _1309_;
  assign _1317_ = _1129_ & _1128_;
  assign _1318_ = ~_1132_;
  assign _temp967_ = _1318_ | _1131_;
  assign _1319_ = ~_temp967_;
  assign _temp968_ = _1319_ | _1317_;
  assign _1320_ = ~_temp968_;
  assign _1321_ = _1320_ ^ _1315_;
  assign _1322_ = ~_1138_;
  assign _temp969_ = _1133_ | _1127_;
  assign _1323_ = ~_temp969_;
  assign _temp970_ = _1322_ & _1134_;
  assign _temp971_ = _temp970_ | _1323_;
  assign _1324_ = ~_temp971_;
  assign _1325_ = _1324_ ^ _1321_;
  assign _temp972_ = b[18] & a[9];
  assign _1326_ = ~_temp972_;
  assign _1328_ = b[19] & a[8];
  assign _1329_ = _1328_ ^ _1326_;
  assign _1330_ = b[20] & a[7];
  assign _1331_ = _1330_ ^ _1329_;
  assign _1332_ = ~_1147_;
  assign _1333_ = _1146_ & _1145_;
  assign _temp973_ = _1148_ & _1332_;
  assign _temp974_ = _temp973_ | _1333_;
  assign _1334_ = ~_temp974_;
  assign _1335_ = _1334_ ^ _1331_;
  assign _1336_ = b[21] & a[6];
  assign _1337_ = b[22] & a[5];
  assign _temp975_ = _1337_ ^ _1336_;
  assign _1339_ = ~_temp975_;
  assign _1340_ = b[23] & a[4];
  assign _1341_ = _1340_ ^ _1339_;
  assign _1342_ = _1341_ ^ _1335_;
  assign _1343_ = _1342_ ^ _1325_;
  assign _1344_ = _1343_ ^ _1306_;
  assign _temp976_ = _1143_ | _1139_;
  assign _1345_ = ~_temp976_;
  assign _1346_ = ~_1160_;
  assign _1347_ = _1346_ & _1144_;
  assign _temp977_ = _1347_ | _1345_;
  assign _1348_ = ~_temp977_;
  assign _1350_ = ~_1348_;
  assign _1351_ = _1350_ ^ _1344_;
  assign _temp978_ = _1351_ ^ _1302_;
  assign _1352_ = ~_temp978_;
  assign _temp979_ = _1120_ | _1116_;
  assign _1353_ = ~_temp979_;
  assign _temp980_ = _1167_ & _1121_;
  assign _temp981_ = _temp980_ | _1353_;
  assign _1354_ = ~_temp981_;
  assign _1355_ = _1354_ ^ _1352_;
  assign _1356_ = _1161_ | _1125_;
  assign _temp982_ = _1166_ | _1162_;
  assign _temp983_ = _temp982_ & _1356_;
  assign _1357_ = ~_temp983_;
  assign _temp984_ = _1151_ | _1149_;
  assign _1358_ = ~_temp984_;
  assign _temp985_ = _1158_ | _1153_;
  assign _1359_ = ~_temp985_;
  assign _temp986_ = _1359_ | _1358_;
  assign _1361_ = ~_temp986_;
  assign _1362_ = ~_1156_;
  assign _1363_ = _1155_ & _1154_;
  assign _temp987_ = _1157_ & _1362_;
  assign _temp988_ = _temp987_ | _1363_;
  assign _1364_ = ~_temp988_;
  assign _temp989_ = b[24] & a[3];
  assign _1365_ = ~_temp989_;
  assign _1366_ = a[2] & b[25];
  assign _1367_ = _1366_ ^ _1365_;
  assign _1368_ = b[26] & a[1];
  assign _1369_ = _1368_ ^ _1367_;
  assign _1370_ = _1369_ ^ _1364_;
  assign _1372_ = _1186_ & _1184_;
  assign _1373_ = ~_1188_;
  assign _temp990_ = _1373_ | _1187_;
  assign _1374_ = ~_temp990_;
  assign _temp991_ = _1374_ | _1372_;
  assign _1375_ = ~_temp991_;
  assign _1376_ = _1375_ ^ _1370_;
  assign _temp992_ = _1376_ ^ _1361_;
  assign _1377_ = ~_temp992_;
  assign _1378_ = ~_1183_;
  assign _temp993_ = _1189_ | _1378_;
  assign _1379_ = ~_temp993_;
  assign _1380_ = ~_1191_;
  assign _temp994_ = _1380_ | _1190_;
  assign _1381_ = ~_temp994_;
  assign _temp995_ = _1381_ | _1379_;
  assign _1383_ = ~_temp995_;
  assign _temp996_ = _1383_ ^ _1377_;
  assign _1384_ = ~_temp996_;
  assign _temp997_ = _1192_ | _1180_;
  assign _1385_ = ~_temp997_;
  assign _temp998_ = _1194_ & _1193_;
  assign _temp999_ = _temp998_ | _1385_;
  assign _1386_ = ~_temp999_;
  assign _temp1000_ = _1386_ ^ _1384_;
  assign _1387_ = ~_temp1000_;
  assign _1388_ = b[27] & a[0];
  assign _1389_ = _1388_ ^ _1387_;
  assign _1390_ = ~_1389_;
  assign _1391_ = _1390_ ^ _1357_;
  assign _temp1001_ = _1199_ | _1195_;
  assign _1392_ = ~_temp1001_;
  assign _1394_ = _1392_ ^ _1391_;
  assign _temp1002_ = _1394_ ^ _1355_;
  assign _1395_ = ~_temp1002_;
  assign _temp1003_ = _1170_ | _1168_;
  assign _1396_ = ~_temp1003_;
  assign _temp1004_ = _1204_ & _1171_;
  assign _temp1005_ = _temp1004_ | _1396_;
  assign _1397_ = ~_temp1005_;
  assign _1398_ = _1397_ ^ _1395_;
  assign _temp1006_ = _1200_ | _1176_;
  assign _1399_ = ~_temp1006_;
  assign _1400_ = _1203_ & _1201_;
  assign _temp1007_ = _1400_ | _1399_;
  assign _1401_ = ~_temp1007_;
  assign _1402_ = _1401_ ^ _1398_;
  assign _temp1008_ = _1208_ | _1205_;
  assign _1403_ = ~_temp1008_;
  assign _temp1009_ = _1212_ & _1209_;
  assign _temp1010_ = _temp1009_ | _1403_;
  assign _1405_ = ~_temp1010_;
  assign _1406_ = _1405_ ^ _1402_;
  assign _temp1011_ = _1215_ | _1213_;
  assign _1407_ = ~_temp1011_;
  assign _1408_ = _1407_ ^ _1406_;
  assign _1409_ = _1217_ & _1216_;
  assign _temp1012_ = _1225_ & _1219_;
  assign _temp1013_ = _temp1012_ | _1409_;
  assign _1410_ = ~_temp1013_;
  assign _temp1014_ = _1410_ ^ _1408_;
  assign q[27] = ~_temp1014_;
  assign _1411_ = a[28] & b[0];
  assign _1412_ = b[1] & a[27];
  assign _temp1015_ = _1412_ ^ _1411_;
  assign _1413_ = ~_temp1015_;
  assign _1415_ = b[2] & a[26];
  assign _1416_ = _1415_ ^ _1413_;
  assign _1417_ = ~_1229_;
  assign _1418_ = _1227_ & _1226_;
  assign _temp1016_ = _1230_ & _1417_;
  assign _temp1017_ = _temp1016_ | _1418_;
  assign _1419_ = ~_temp1017_;
  assign _temp1018_ = _1419_ ^ _1416_;
  assign _1420_ = ~_temp1018_;
  assign _1421_ = b[3] & a[25];
  assign _1422_ = b[4] & a[24];
  assign _temp1019_ = _1422_ ^ _1421_;
  assign _1423_ = ~_temp1019_;
  assign _1424_ = b[5] & a[23];
  assign _1426_ = _1424_ ^ _1423_;
  assign _1427_ = ~_1426_;
  assign _1428_ = _1427_ ^ _1420_;
  assign _temp1020_ = _1233_ | _1231_;
  assign _1429_ = ~_temp1020_;
  assign _temp1021_ = _1240_ | _1234_;
  assign _1430_ = ~_temp1021_;
  assign _temp1022_ = _1430_ | _1429_;
  assign _1431_ = ~_temp1022_;
  assign _temp1023_ = _1431_ ^ _1428_;
  assign _1432_ = ~_temp1023_;
  assign _1433_ = ~_1235_;
  assign _1434_ = _1236_ & _1433_;
  assign _1435_ = ~_1238_;
  assign _temp1024_ = _1435_ | _1237_;
  assign _1436_ = ~_temp1024_;
  assign _temp1025_ = _1436_ | _1434_;
  assign _1437_ = ~_temp1025_;
  assign _1438_ = b[6] & a[22];
  assign _1439_ = b[7] & a[21];
  assign _temp1026_ = _1439_ ^ _1438_;
  assign _1440_ = ~_temp1026_;
  assign _1441_ = b[8] & a[20];
  assign _1442_ = _1441_ ^ _1440_;
  assign _temp1027_ = _1442_ ^ _1437_;
  assign _1443_ = ~_temp1027_;
  assign _1444_ = ~_1252_;
  assign _1445_ = _1253_ & _1444_;
  assign _1447_ = ~_1255_;
  assign _temp1028_ = _1447_ | _1254_;
  assign _1448_ = ~_temp1028_;
  assign _temp1029_ = _1448_ | _1445_;
  assign _1449_ = ~_temp1029_;
  assign _1450_ = ~_1449_;
  assign _1451_ = _1450_ ^ _1443_;
  assign _1452_ = ~_1451_;
  assign _1453_ = _1452_ ^ _1432_;
  assign _temp1030_ = _1245_ | _1242_;
  assign _1454_ = ~_temp1030_;
  assign _temp1031_ = _1264_ | _1246_;
  assign _1455_ = ~_temp1031_;
  assign _temp1032_ = _1455_ | _1454_;
  assign _1456_ = ~_temp1032_;
  assign _temp1033_ = _1456_ ^ _1453_;
  assign _1458_ = ~_temp1033_;
  assign _temp1034_ = _1256_ | _1251_;
  assign _1459_ = ~_temp1034_;
  assign _temp1035_ = _1262_ | _1257_;
  assign _1460_ = ~_temp1035_;
  assign _temp1036_ = _1460_ | _1459_;
  assign _1461_ = ~_temp1036_;
  assign _1462_ = b[9] & a[19];
  assign _1463_ = b[10] & a[18];
  assign _temp1037_ = _1463_ ^ _1462_;
  assign _1464_ = ~_temp1037_;
  assign _1465_ = b[11] & a[17];
  assign _1466_ = _1465_ ^ _1464_;
  assign _1467_ = ~_1277_;
  assign _1469_ = ~_1275_;
  assign _1470_ = _1276_ & _1469_;
  assign _temp1038_ = _1278_ & _1467_;
  assign _temp1039_ = _temp1038_ | _1470_;
  assign _1471_ = ~_temp1039_;
  assign _1472_ = _1471_ ^ _1466_;
  assign _1473_ = b[12] & a[16];
  assign _1474_ = b[13] & a[15];
  assign _temp1040_ = _1474_ ^ _1473_;
  assign _1475_ = ~_temp1040_;
  assign _1476_ = b[14] & a[14];
  assign _1477_ = _1476_ ^ _1475_;
  assign _1478_ = _1477_ ^ _1472_;
  assign _temp1041_ = _1478_ ^ _1461_;
  assign _1480_ = ~_temp1041_;
  assign _temp1042_ = _1282_ | _1279_;
  assign _1481_ = ~_temp1042_;
  assign _1482_ = ~_1289_;
  assign _1483_ = _1482_ & _1284_;
  assign _temp1043_ = _1483_ | _1481_;
  assign _1484_ = ~_temp1043_;
  assign _1485_ = ~_1484_;
  assign _1486_ = _1485_ ^ _1480_;
  assign _temp1044_ = _1486_ ^ _1458_;
  assign _1487_ = ~_temp1044_;
  assign _temp1045_ = _1268_ | _1265_;
  assign _1488_ = ~_temp1045_;
  assign _temp1046_ = _1298_ & _1269_;
  assign _temp1047_ = _temp1046_ | _1488_;
  assign _1489_ = ~_temp1047_;
  assign _temp1048_ = _1489_ ^ _1487_;
  assign _1491_ = ~_temp1048_;
  assign _1492_ = ~_1491_;
  assign _temp1049_ = _1290_ | _1274_;
  assign _1493_ = ~_temp1049_;
  assign _1494_ = _1297_ & _1291_;
  assign _temp1050_ = _1494_ | _1493_;
  assign _1495_ = ~_temp1050_;
  assign _1496_ = ~_1287_;
  assign _1497_ = ~_1285_;
  assign _1498_ = _1286_ & _1497_;
  assign _temp1051_ = _1288_ & _1496_;
  assign _temp1052_ = _temp1051_ | _1498_;
  assign _1499_ = ~_temp1052_;
  assign _1500_ = b[15] & a[13];
  assign _1502_ = b[16] & a[12];
  assign _temp1053_ = _1502_ ^ _1500_;
  assign _1503_ = ~_temp1053_;
  assign _1504_ = b[17] & a[11];
  assign _1505_ = _1504_ ^ _1503_;
  assign _1506_ = _1505_ ^ _1499_;
  assign _1507_ = ~_1310_;
  assign _1508_ = _1311_ & _1507_;
  assign _1509_ = ~_1313_;
  assign _temp1054_ = _1509_ | _1312_;
  assign _1510_ = ~_temp1054_;
  assign _temp1055_ = _1510_ | _1508_;
  assign _1511_ = ~_temp1055_;
  assign _1513_ = _1511_ ^ _1506_;
  assign _1514_ = ~_1320_;
  assign _temp1056_ = _1314_ | _1309_;
  assign _1515_ = ~_temp1056_;
  assign _temp1057_ = _1514_ & _1315_;
  assign _temp1058_ = _temp1057_ | _1515_;
  assign _1516_ = ~_temp1058_;
  assign _1517_ = _1516_ ^ _1513_;
  assign _1518_ = b[18] & a[10];
  assign _1519_ = b[19] & a[9];
  assign _temp1059_ = _1519_ ^ _1518_;
  assign _1520_ = ~_temp1059_;
  assign _1521_ = b[20] & a[8];
  assign _1522_ = _1521_ ^ _1520_;
  assign _1524_ = ~_1329_;
  assign _1525_ = ~_1326_;
  assign _1526_ = _1328_ & _1525_;
  assign _temp1060_ = _1330_ & _1524_;
  assign _temp1061_ = _temp1060_ | _1526_;
  assign _1527_ = ~_temp1061_;
  assign _1528_ = _1527_ ^ _1522_;
  assign _1529_ = b[21] & a[7];
  assign _1530_ = b[22] & a[6];
  assign _temp1062_ = _1530_ ^ _1529_;
  assign _1531_ = ~_temp1062_;
  assign _1532_ = b[23] & a[5];
  assign _1533_ = _1532_ ^ _1531_;
  assign _1535_ = _1533_ ^ _1528_;
  assign _1536_ = _1535_ ^ _1517_;
  assign _1537_ = _1536_ ^ _1495_;
  assign _temp1063_ = _1324_ | _1321_;
  assign _1538_ = ~_temp1063_;
  assign _1539_ = ~_1342_;
  assign _1540_ = _1539_ & _1325_;
  assign _temp1064_ = _1540_ | _1538_;
  assign _1541_ = ~_temp1064_;
  assign _1542_ = _1541_ ^ _1537_;
  assign _1543_ = _1542_ ^ _1492_;
  assign _temp1065_ = _1301_ | _1299_;
  assign _1544_ = ~_temp1065_;
  assign _temp1066_ = _1351_ & _1302_;
  assign _temp1067_ = _temp1066_ | _1544_;
  assign _1546_ = ~_temp1067_;
  assign _1547_ = _1546_ ^ _1543_;
  assign _temp1068_ = _1343_ | _1306_;
  assign _1548_ = ~_temp1068_;
  assign _1549_ = _1350_ & _1344_;
  assign _temp1069_ = _1549_ | _1548_;
  assign _1550_ = ~_temp1069_;
  assign _1551_ = ~_1341_;
  assign _temp1070_ = _1334_ | _1331_;
  assign _1552_ = ~_temp1070_;
  assign _temp1071_ = _1551_ & _1335_;
  assign _temp1072_ = _temp1071_ | _1552_;
  assign _1553_ = ~_temp1072_;
  assign _1554_ = ~_1339_;
  assign _1555_ = _1337_ & _1336_;
  assign _temp1073_ = _1340_ & _1554_;
  assign _temp1074_ = _temp1073_ | _1555_;
  assign _1557_ = ~_temp1074_;
  assign _1558_ = a[4] & b[24];
  assign _1559_ = b[25] & a[3];
  assign _temp1075_ = _1559_ ^ _1558_;
  assign _1560_ = ~_temp1075_;
  assign _1561_ = b[26] & a[2];
  assign _1562_ = _1561_ ^ _1560_;
  assign _1563_ = _1562_ ^ _1557_;
  assign _1564_ = ~_1365_;
  assign _1565_ = _1366_ & _1564_;
  assign _1566_ = ~_1368_;
  assign _temp1076_ = _1566_ | _1367_;
  assign _1568_ = ~_temp1076_;
  assign _temp1077_ = _1568_ | _1565_;
  assign _1569_ = ~_temp1077_;
  assign _1570_ = _1569_ ^ _1563_;
  assign _1571_ = _1570_ ^ _1553_;
  assign _temp1078_ = _1369_ | _1364_;
  assign _1572_ = ~_temp1078_;
  assign _1573_ = ~_1375_;
  assign _1574_ = _1573_ & _1370_;
  assign _temp1079_ = _1574_ | _1572_;
  assign _1575_ = ~_temp1079_;
  assign _1576_ = _1575_ ^ _1571_;
  assign _temp1080_ = _1376_ | _1361_;
  assign _1577_ = ~_temp1080_;
  assign _temp1081_ = _1383_ | _1377_;
  assign _1579_ = ~_temp1081_;
  assign _temp1082_ = _1579_ | _1577_;
  assign _1580_ = ~_temp1082_;
  assign _1581_ = _1580_ ^ _1576_;
  assign _1582_ = b[27] & a[1];
  assign _1583_ = b[28] & a[0];
  assign _temp1083_ = _1583_ ^ _1582_;
  assign _1584_ = ~_temp1083_;
  assign _1585_ = _1584_ ^ _1581_;
  assign _1586_ = _1585_ ^ _1550_;
  assign _temp1084_ = _1386_ | _1384_;
  assign _1587_ = ~_temp1084_;
  assign _1588_ = ~_1388_;
  assign _temp1085_ = _1588_ | _1387_;
  assign _1590_ = ~_temp1085_;
  assign _temp1086_ = _1590_ | _1587_;
  assign _1591_ = ~_temp1086_;
  assign _1592_ = ~_1591_;
  assign _1593_ = _1592_ ^ _1586_;
  assign _temp1087_ = _1593_ ^ _1547_;
  assign _1594_ = ~_temp1087_;
  assign _temp1088_ = _1354_ | _1352_;
  assign _1595_ = ~_temp1088_;
  assign _temp1089_ = _1394_ & _1355_;
  assign _temp1090_ = _temp1089_ | _1595_;
  assign _1596_ = ~_temp1090_;
  assign _1597_ = _1596_ ^ _1594_;
  assign _1598_ = _1390_ & _1357_;
  assign _1599_ = _1392_ & _1391_;
  assign _temp1091_ = _1599_ | _1598_;
  assign _1601_ = ~_temp1091_;
  assign _1602_ = _1601_ ^ _1597_;
  assign _1603_ = ~_1401_;
  assign _temp1092_ = _1397_ | _1395_;
  assign _1604_ = ~_temp1092_;
  assign _temp1093_ = _1603_ & _1398_;
  assign _temp1094_ = _temp1093_ | _1604_;
  assign _1605_ = ~_temp1094_;
  assign _1606_ = _1605_ ^ _1602_;
  assign _temp1095_ = _1405_ | _1402_;
  assign _1607_ = ~_temp1095_;
  assign _temp1096_ = _1607_ ^ _1606_;
  assign _1608_ = ~_temp1096_;
  assign _temp1097_ = _1408_ & _1219_;
  assign _1609_ = ~_temp1097_;
  assign _temp1098_ = _1609_ | _1224_;
  assign _1610_ = ~_temp1098_;
  assign _1612_ = _1407_ & _1406_;
  assign _temp1099_ = _1409_ & _1408_;
  assign _temp1100_ = _temp1099_ | _1612_;
  assign _1613_ = ~_temp1100_;
  assign _temp1101_ = _1609_ | _1223_;
  assign _temp1102_ = _temp1101_ & _1613_;
  assign _1614_ = ~_temp1102_;
  assign _temp1103_ = _1610_ & _0887_;
  assign _temp1104_ = _temp1103_ | _1614_;
  assign _1615_ = ~_temp1104_;
  assign q[28] = _1615_ ^ _1608_;
  assign _1616_ = a[29] & b[0];
  assign _1617_ = b[1] & a[28];
  assign _temp1105_ = _1617_ ^ _1616_;
  assign _1618_ = ~_temp1105_;
  assign _1619_ = b[2] & a[27];
  assign _1620_ = _1619_ ^ _1618_;
  assign _1622_ = ~_1413_;
  assign _1623_ = _1412_ & _1411_;
  assign _temp1106_ = _1415_ & _1622_;
  assign _temp1107_ = _temp1106_ | _1623_;
  assign _1624_ = ~_temp1107_;
  assign _temp1108_ = _1624_ ^ _1620_;
  assign _1625_ = ~_temp1108_;
  assign _1626_ = b[3] & a[26];
  assign _1627_ = b[4] & a[25];
  assign _temp1109_ = _1627_ ^ _1626_;
  assign _1628_ = ~_temp1109_;
  assign _1629_ = b[5] & a[24];
  assign _1630_ = _1629_ ^ _1628_;
  assign _1631_ = ~_1630_;
  assign _1633_ = _1631_ ^ _1625_;
  assign _temp1110_ = _1419_ | _1416_;
  assign _1634_ = ~_temp1110_;
  assign _temp1111_ = _1426_ | _1420_;
  assign _1635_ = ~_temp1111_;
  assign _temp1112_ = _1635_ | _1634_;
  assign _1636_ = ~_temp1112_;
  assign _temp1113_ = _1636_ ^ _1633_;
  assign _1637_ = ~_temp1113_;
  assign _1638_ = ~_1423_;
  assign _1639_ = _1422_ & _1421_;
  assign _temp1114_ = _1424_ & _1638_;
  assign _temp1115_ = _temp1114_ | _1639_;
  assign _1640_ = ~_temp1115_;
  assign _1641_ = b[6] & a[23];
  assign _1642_ = b[7] & a[22];
  assign _temp1116_ = _1642_ ^ _1641_;
  assign _1644_ = ~_temp1116_;
  assign _1645_ = b[8] & a[21];
  assign _1646_ = _1645_ ^ _1644_;
  assign _1647_ = _1646_ ^ _1640_;
  assign _1648_ = _1439_ & _1438_;
  assign _1649_ = ~_1441_;
  assign _temp1117_ = _1649_ | _1440_;
  assign _1650_ = ~_temp1117_;
  assign _temp1118_ = _1650_ | _1648_;
  assign _1651_ = ~_temp1118_;
  assign _1652_ = _1651_ ^ _1647_;
  assign _1653_ = ~_1652_;
  assign _1655_ = _1653_ ^ _1637_;
  assign _temp1119_ = _1431_ | _1428_;
  assign _1656_ = ~_temp1119_;
  assign _temp1120_ = _1451_ | _1432_;
  assign _1657_ = ~_temp1120_;
  assign _temp1121_ = _1657_ | _1656_;
  assign _1658_ = ~_temp1121_;
  assign _temp1122_ = _1658_ ^ _1655_;
  assign _1659_ = ~_temp1122_;
  assign _temp1123_ = _1442_ | _1437_;
  assign _1660_ = ~_temp1123_;
  assign _temp1124_ = _1449_ | _1443_;
  assign _1661_ = ~_temp1124_;
  assign _temp1125_ = _1661_ | _1660_;
  assign _1662_ = ~_temp1125_;
  assign _1663_ = b[9] & a[20];
  assign _1664_ = b[10] & a[19];
  assign _temp1126_ = _1664_ ^ _1663_;
  assign _1666_ = ~_temp1126_;
  assign _1667_ = b[11] & a[18];
  assign _1668_ = _1667_ ^ _1666_;
  assign _1669_ = ~_1464_;
  assign _1670_ = _1463_ & _1462_;
  assign _temp1127_ = _1465_ & _1669_;
  assign _temp1128_ = _temp1127_ | _1670_;
  assign _1671_ = ~_temp1128_;
  assign _1672_ = _1671_ ^ _1668_;
  assign _1673_ = b[12] & a[17];
  assign _1674_ = b[13] & a[16];
  assign _temp1129_ = _1674_ ^ _1673_;
  assign _1675_ = ~_temp1129_;
  assign _1677_ = b[14] & a[15];
  assign _1678_ = _1677_ ^ _1675_;
  assign _1679_ = _1678_ ^ _1672_;
  assign _1680_ = _1679_ ^ _1662_;
  assign _temp1130_ = _1471_ | _1466_;
  assign _1681_ = ~_temp1130_;
  assign _1682_ = ~_1477_;
  assign _1683_ = _1682_ & _1472_;
  assign _temp1131_ = _1683_ | _1681_;
  assign _1684_ = ~_temp1131_;
  assign _1685_ = _1684_ ^ _1680_;
  assign _1686_ = ~_1685_;
  assign _1688_ = _1686_ ^ _1659_;
  assign _temp1132_ = _1456_ | _1453_;
  assign _1689_ = ~_temp1132_;
  assign _temp1133_ = _1486_ | _1458_;
  assign _1690_ = ~_temp1133_;
  assign _temp1134_ = _1690_ | _1689_;
  assign _1691_ = ~_temp1134_;
  assign _temp1135_ = _1691_ ^ _1688_;
  assign _1692_ = ~_temp1135_;
  assign _temp1136_ = _1478_ | _1461_;
  assign _1693_ = ~_temp1136_;
  assign _temp1137_ = _1484_ | _1480_;
  assign _1694_ = ~_temp1137_;
  assign _temp1138_ = _1694_ | _1693_;
  assign _1695_ = ~_temp1138_;
  assign _1696_ = ~_1475_;
  assign _1697_ = _1474_ & _1473_;
  assign _temp1139_ = _1476_ & _1696_;
  assign _temp1140_ = _temp1139_ | _1697_;
  assign _1699_ = ~_temp1140_;
  assign _1700_ = b[15] & a[14];
  assign _1701_ = b[16] & a[13];
  assign _temp1141_ = _1701_ ^ _1700_;
  assign _1702_ = ~_temp1141_;
  assign _1703_ = b[17] & a[12];
  assign _1704_ = _1703_ ^ _1702_;
  assign _1705_ = _1704_ ^ _1699_;
  assign _1706_ = _1502_ & _1500_;
  assign _1707_ = ~_1504_;
  assign _temp1142_ = _1707_ | _1503_;
  assign _1708_ = ~_temp1142_;
  assign _temp1143_ = _1708_ | _1706_;
  assign _1710_ = ~_temp1143_;
  assign _1711_ = _1710_ ^ _1705_;
  assign _1712_ = ~_1511_;
  assign _temp1144_ = _1505_ | _1499_;
  assign _1713_ = ~_temp1144_;
  assign _temp1145_ = _1712_ & _1506_;
  assign _temp1146_ = _temp1145_ | _1713_;
  assign _1714_ = ~_temp1146_;
  assign _1715_ = _1714_ ^ _1711_;
  assign _1716_ = b[18] & a[11];
  assign _1717_ = b[19] & a[10];
  assign _temp1147_ = _1717_ ^ _1716_;
  assign _1718_ = ~_temp1147_;
  assign _1719_ = b[20] & a[9];
  assign _1721_ = _1719_ ^ _1718_;
  assign _1722_ = ~_1520_;
  assign _1723_ = _1519_ & _1518_;
  assign _temp1148_ = _1521_ & _1722_;
  assign _temp1149_ = _temp1148_ | _1723_;
  assign _1724_ = ~_temp1149_;
  assign _temp1150_ = _1724_ ^ _1721_;
  assign _1725_ = ~_temp1150_;
  assign _1726_ = b[21] & a[8];
  assign _1727_ = b[22] & a[7];
  assign _temp1151_ = _1727_ ^ _1726_;
  assign _1728_ = ~_temp1151_;
  assign _1729_ = b[23] & a[6];
  assign _1730_ = _1729_ ^ _1728_;
  assign _1732_ = ~_1730_;
  assign _1733_ = _1732_ ^ _1725_;
  assign _1734_ = _1733_ ^ _1715_;
  assign _temp1152_ = _1734_ ^ _1695_;
  assign _1735_ = ~_temp1152_;
  assign _temp1153_ = _1516_ | _1513_;
  assign _1736_ = ~_temp1153_;
  assign _1737_ = ~_1535_;
  assign _1738_ = _1737_ & _1517_;
  assign _temp1154_ = _1738_ | _1736_;
  assign _1739_ = ~_temp1154_;
  assign _1740_ = ~_1739_;
  assign _1741_ = _1740_ ^ _1735_;
  assign _temp1155_ = _1741_ ^ _1692_;
  assign _1743_ = ~_temp1155_;
  assign _temp1156_ = _1489_ | _1487_;
  assign _1744_ = ~_temp1156_;
  assign _temp1157_ = _1542_ | _1491_;
  assign _1745_ = ~_temp1157_;
  assign _temp1158_ = _1745_ | _1744_;
  assign _1746_ = ~_temp1158_;
  assign _temp1159_ = _1746_ ^ _1743_;
  assign _1747_ = ~_temp1159_;
  assign _temp1160_ = _1536_ | _1495_;
  assign _1748_ = ~_temp1160_;
  assign _1749_ = ~_1541_;
  assign _1750_ = _1749_ & _1537_;
  assign _temp1161_ = _1750_ | _1748_;
  assign _1751_ = ~_temp1161_;
  assign _1752_ = ~_1533_;
  assign _temp1162_ = _1527_ | _1522_;
  assign _1754_ = ~_temp1162_;
  assign _temp1163_ = _1752_ & _1528_;
  assign _temp1164_ = _temp1163_ | _1754_;
  assign _1755_ = ~_temp1164_;
  assign _1756_ = ~_1531_;
  assign _1757_ = _1530_ & _1529_;
  assign _temp1165_ = _1532_ & _1756_;
  assign _temp1166_ = _temp1165_ | _1757_;
  assign _1758_ = ~_temp1166_;
  assign _1759_ = a[5] & b[24];
  assign _1760_ = b[25] & a[4];
  assign _temp1167_ = _1760_ ^ _1759_;
  assign _1761_ = ~_temp1167_;
  assign _1762_ = b[26] & a[3];
  assign _1763_ = _1762_ ^ _1761_;
  assign _1765_ = _1763_ ^ _1758_;
  assign _1766_ = _1559_ & _1558_;
  assign _1767_ = ~_1561_;
  assign _temp1168_ = _1767_ | _1560_;
  assign _1768_ = ~_temp1168_;
  assign _temp1169_ = _1768_ | _1766_;
  assign _1769_ = ~_temp1169_;
  assign _1770_ = _1769_ ^ _1765_;
  assign _1771_ = _1770_ ^ _1755_;
  assign _temp1170_ = _1562_ | _1557_;
  assign _1772_ = ~_temp1170_;
  assign _1773_ = ~_1569_;
  assign _1774_ = _1773_ & _1563_;
  assign _temp1171_ = _1774_ | _1772_;
  assign _1776_ = ~_temp1171_;
  assign _1777_ = _1776_ ^ _1771_;
  assign _1778_ = ~_1575_;
  assign _temp1172_ = _1570_ | _1553_;
  assign _1779_ = ~_temp1172_;
  assign _temp1173_ = _1778_ & _1571_;
  assign _temp1174_ = _temp1173_ | _1779_;
  assign _1780_ = ~_temp1174_;
  assign _1781_ = _1780_ ^ _1777_;
  assign _1782_ = b[27] & a[2];
  assign _1783_ = b[28] & a[1];
  assign _temp1175_ = _1783_ ^ _1782_;
  assign _1784_ = ~_temp1175_;
  assign _1785_ = b[29] & a[0];
  assign _1787_ = _1785_ ^ _1784_;
  assign _1788_ = _1583_ & _1582_;
  assign _1789_ = _1788_ ^ _1787_;
  assign _1790_ = _1789_ ^ _1781_;
  assign _1791_ = _1790_ ^ _1751_;
  assign _temp1176_ = _1580_ | _1576_;
  assign _1792_ = ~_temp1176_;
  assign _1793_ = ~_1584_;
  assign _1794_ = _1793_ & _1581_;
  assign _temp1177_ = _1794_ | _1792_;
  assign _1795_ = ~_temp1177_;
  assign _1796_ = _1795_ ^ _1791_;
  assign _1798_ = _1796_ ^ _1747_;
  assign _temp1178_ = _1546_ | _1543_;
  assign _1799_ = ~_temp1178_;
  assign _temp1179_ = _1593_ & _1547_;
  assign _temp1180_ = _temp1179_ | _1799_;
  assign _1800_ = ~_temp1180_;
  assign _1801_ = _1800_ ^ _1798_;
  assign _temp1181_ = _1585_ | _1550_;
  assign _1802_ = ~_temp1181_;
  assign _1803_ = _1592_ & _1586_;
  assign _temp1182_ = _1803_ | _1802_;
  assign _1804_ = ~_temp1182_;
  assign _1805_ = _1804_ ^ _1801_;
  assign _1806_ = ~_1601_;
  assign _temp1183_ = _1806_ & _1597_;
  assign _1807_ = ~_temp1183_;
  assign _temp1184_ = _1596_ | _1594_;
  assign _temp1185_ = _temp1184_ & _1807_;
  assign _1809_ = ~_temp1185_;
  assign _1810_ = _1809_ ^ _1805_;
  assign _temp1186_ = _1605_ | _1602_;
  assign _1811_ = ~_temp1186_;
  assign _1812_ = _1811_ ^ _1810_;
  assign _1813_ = _1607_ & _1606_;
  assign _1814_ = ~_1813_;
  assign _temp1187_ = _1615_ | _1608_;
  assign _temp1188_ = _temp1187_ & _1814_;
  assign _1815_ = ~_temp1188_;
  assign q[29] = _1815_ ^ _1812_;
  assign _1816_ = a[30] & b[0];
  assign _1817_ = b[1] & a[29];
  assign _temp1189_ = _1817_ ^ _1816_;
  assign _1819_ = ~_temp1189_;
  assign _1820_ = b[2] & a[28];
  assign _1821_ = _1820_ ^ _1819_;
  assign _1822_ = ~_1618_;
  assign _1823_ = _1617_ & _1616_;
  assign _temp1190_ = _1619_ & _1822_;
  assign _temp1191_ = _temp1190_ | _1823_;
  assign _1824_ = ~_temp1191_;
  assign _temp1192_ = _1824_ ^ _1821_;
  assign _1825_ = ~_temp1192_;
  assign _1826_ = b[3] & a[27];
  assign _1827_ = b[4] & a[26];
  assign _temp1193_ = _1827_ ^ _1826_;
  assign _1828_ = ~_temp1193_;
  assign _1830_ = b[5] & a[25];
  assign _1831_ = _1830_ ^ _1828_;
  assign _temp1194_ = _1831_ ^ _1825_;
  assign _1832_ = ~_temp1194_;
  assign _temp1195_ = _1624_ | _1620_;
  assign _1833_ = ~_temp1195_;
  assign _temp1196_ = _1630_ | _1625_;
  assign _1834_ = ~_temp1196_;
  assign _temp1197_ = _1834_ | _1833_;
  assign _1835_ = ~_temp1197_;
  assign _1836_ = _1835_ ^ _1832_;
  assign _1837_ = ~_1628_;
  assign _1838_ = _1627_ & _1626_;
  assign _temp1198_ = _1629_ & _1837_;
  assign _temp1199_ = _temp1198_ | _1838_;
  assign _1839_ = ~_temp1199_;
  assign _1841_ = b[6] & a[24];
  assign _1842_ = b[7] & a[23];
  assign _temp1200_ = _1842_ ^ _1841_;
  assign _1843_ = ~_temp1200_;
  assign _1844_ = b[8] & a[22];
  assign _1845_ = _1844_ ^ _1843_;
  assign _temp1201_ = _1845_ ^ _1839_;
  assign _1846_ = ~_temp1201_;
  assign _1847_ = _1642_ & _1641_;
  assign _1848_ = ~_1645_;
  assign _temp1202_ = _1848_ | _1644_;
  assign _1849_ = ~_temp1202_;
  assign _temp1203_ = _1849_ | _1847_;
  assign _1850_ = ~_temp1203_;
  assign _temp1204_ = _1850_ ^ _1846_;
  assign _1852_ = ~_temp1204_;
  assign _1853_ = ~_1852_;
  assign _1854_ = _1853_ ^ _1836_;
  assign _1855_ = _1636_ | _1633_;
  assign _temp1205_ = _1652_ | _1637_;
  assign _temp1206_ = _temp1205_ & _1855_;
  assign _1856_ = ~_temp1206_;
  assign _1857_ = _1856_ ^ _1854_;
  assign _1858_ = ~_1651_;
  assign _temp1207_ = _1646_ | _1640_;
  assign _1859_ = ~_temp1207_;
  assign _temp1208_ = _1858_ & _1647_;
  assign _temp1209_ = _temp1208_ | _1859_;
  assign _1860_ = ~_temp1209_;
  assign _1861_ = b[9] & a[21];
  assign _1863_ = b[10] & a[20];
  assign _temp1210_ = _1863_ ^ _1861_;
  assign _1864_ = ~_temp1210_;
  assign _1865_ = b[11] & a[19];
  assign _1866_ = _1865_ ^ _1864_;
  assign _1867_ = ~_1666_;
  assign _1868_ = _1664_ & _1663_;
  assign _temp1211_ = _1667_ & _1867_;
  assign _temp1212_ = _temp1211_ | _1868_;
  assign _1869_ = ~_temp1212_;
  assign _temp1213_ = _1869_ ^ _1866_;
  assign _1870_ = ~_temp1213_;
  assign _1871_ = b[12] & a[18];
  assign _1872_ = b[13] & a[17];
  assign _temp1214_ = _1872_ ^ _1871_;
  assign _1874_ = ~_temp1214_;
  assign _1875_ = b[14] & a[16];
  assign _1876_ = _1875_ ^ _1874_;
  assign _1877_ = ~_1876_;
  assign _1878_ = _1877_ ^ _1870_;
  assign _temp1215_ = _1878_ ^ _1860_;
  assign _1879_ = ~_temp1215_;
  assign _temp1216_ = _1671_ | _1668_;
  assign _1880_ = ~_temp1216_;
  assign _1881_ = ~_1678_;
  assign _1882_ = _1881_ & _1672_;
  assign _temp1217_ = _1882_ | _1880_;
  assign _1883_ = ~_temp1217_;
  assign _temp1218_ = _1883_ ^ _1879_;
  assign _1885_ = ~_temp1218_;
  assign _1886_ = ~_1885_;
  assign _1887_ = _1886_ ^ _1857_;
  assign _1888_ = _1658_ | _1655_;
  assign _temp1219_ = _1685_ | _1659_;
  assign _temp1220_ = _temp1219_ & _1888_;
  assign _1889_ = ~_temp1220_;
  assign _1890_ = _1889_ ^ _1887_;
  assign _1891_ = ~_1684_;
  assign _temp1221_ = _1891_ & _1680_;
  assign _1892_ = ~_temp1221_;
  assign _temp1222_ = _1679_ | _1662_;
  assign _temp1223_ = _temp1222_ & _1892_;
  assign _1893_ = ~_temp1223_;
  assign _1894_ = ~_1675_;
  assign _1896_ = _1674_ & _1673_;
  assign _temp1224_ = _1677_ & _1894_;
  assign _temp1225_ = _temp1224_ | _1896_;
  assign _1897_ = ~_temp1225_;
  assign _1898_ = b[15] & a[15];
  assign _1899_ = b[16] & a[14];
  assign _temp1226_ = _1899_ ^ _1898_;
  assign _1900_ = ~_temp1226_;
  assign _1901_ = b[17] & a[13];
  assign _1902_ = _1901_ ^ _1900_;
  assign _temp1227_ = _1902_ ^ _1897_;
  assign _1903_ = ~_temp1227_;
  assign _1904_ = _1701_ & _1700_;
  assign _1905_ = ~_1703_;
  assign _temp1228_ = _1905_ | _1702_;
  assign _1906_ = ~_temp1228_;
  assign _temp1229_ = _1906_ | _1904_;
  assign _1907_ = ~_temp1229_;
  assign _1908_ = ~_1907_;
  assign _1909_ = _1908_ ^ _1903_;
  assign _1910_ = ~_1710_;
  assign _temp1230_ = _1704_ | _1699_;
  assign _1911_ = ~_temp1230_;
  assign _temp1231_ = _1910_ & _1705_;
  assign _temp1232_ = _temp1231_ | _1911_;
  assign _1912_ = ~_temp1232_;
  assign _temp1233_ = _1912_ ^ _1909_;
  assign _1913_ = ~_temp1233_;
  assign _1914_ = b[18] & a[12];
  assign _1915_ = b[19] & a[11];
  assign _temp1234_ = _1915_ ^ _1914_;
  assign _1917_ = ~_temp1234_;
  assign _1918_ = b[20] & a[10];
  assign _1919_ = _1918_ ^ _1917_;
  assign _1920_ = ~_1718_;
  assign _1921_ = _1717_ & _1716_;
  assign _temp1235_ = _1719_ & _1920_;
  assign _temp1236_ = _temp1235_ | _1921_;
  assign _1922_ = ~_temp1236_;
  assign _temp1237_ = _1922_ ^ _1919_;
  assign _1923_ = ~_temp1237_;
  assign _1924_ = b[21] & a[9];
  assign _1925_ = b[22] & a[8];
  assign _temp1238_ = _1925_ ^ _1924_;
  assign _1926_ = ~_temp1238_;
  assign _1928_ = b[23] & a[7];
  assign _1929_ = _1928_ ^ _1926_;
  assign _1930_ = ~_1929_;
  assign _1931_ = _1930_ ^ _1923_;
  assign _temp1239_ = _1931_ ^ _1913_;
  assign _1932_ = ~_temp1239_;
  assign _1933_ = ~_1932_;
  assign _1934_ = _1933_ ^ _1893_;
  assign _1935_ = ~_1733_;
  assign _temp1240_ = _1714_ | _1711_;
  assign _1936_ = ~_temp1240_;
  assign _temp1241_ = _1935_ & _1715_;
  assign _temp1242_ = _temp1241_ | _1936_;
  assign _1937_ = ~_temp1242_;
  assign _1939_ = ~_1937_;
  assign _1940_ = _1939_ ^ _1934_;
  assign _1941_ = _1940_ ^ _1890_;
  assign _1942_ = _1691_ | _1688_;
  assign _temp1243_ = _1741_ | _1692_;
  assign _temp1244_ = _temp1243_ & _1942_;
  assign _1943_ = ~_temp1244_;
  assign _1944_ = _1943_ ^ _1941_;
  assign _1945_ = _1734_ | _1695_;
  assign _temp1245_ = _1739_ | _1735_;
  assign _temp1246_ = _temp1245_ & _1945_;
  assign _1946_ = ~_temp1246_;
  assign _temp1247_ = _1724_ | _1721_;
  assign _1947_ = ~_temp1247_;
  assign _temp1248_ = _1730_ | _1725_;
  assign _1948_ = ~_temp1248_;
  assign _temp1249_ = _1948_ | _1947_;
  assign _1950_ = ~_temp1249_;
  assign _1951_ = ~_1728_;
  assign _1952_ = _1727_ & _1726_;
  assign _temp1250_ = _1729_ & _1951_;
  assign _temp1251_ = _temp1250_ | _1952_;
  assign _1953_ = ~_temp1251_;
  assign _1954_ = a[6] & b[24];
  assign _1955_ = b[25] & a[5];
  assign _temp1252_ = _1955_ ^ _1954_;
  assign _1956_ = ~_temp1252_;
  assign _1957_ = b[26] & a[4];
  assign _1958_ = _1957_ ^ _1956_;
  assign _temp1253_ = _1958_ ^ _1953_;
  assign _1959_ = ~_temp1253_;
  assign _1961_ = _1760_ & _1759_;
  assign _1962_ = ~_1762_;
  assign _temp1254_ = _1962_ | _1761_;
  assign _1963_ = ~_temp1254_;
  assign _temp1255_ = _1963_ | _1961_;
  assign _1964_ = ~_temp1255_;
  assign _1965_ = ~_1964_;
  assign _1966_ = _1965_ ^ _1959_;
  assign _temp1256_ = _1966_ ^ _1950_;
  assign _1967_ = ~_temp1256_;
  assign _temp1257_ = _1763_ | _1758_;
  assign _1968_ = ~_temp1257_;
  assign _1969_ = ~_1769_;
  assign _1970_ = _1969_ & _1765_;
  assign _temp1258_ = _1970_ | _1968_;
  assign _1972_ = ~_temp1258_;
  assign _temp1259_ = _1972_ ^ _1967_;
  assign _1973_ = ~_temp1259_;
  assign _1974_ = ~_1776_;
  assign _temp1260_ = _1770_ | _1755_;
  assign _1975_ = ~_temp1260_;
  assign _temp1261_ = _1974_ & _1771_;
  assign _temp1262_ = _temp1261_ | _1975_;
  assign _1976_ = ~_temp1262_;
  assign _1977_ = _1976_ ^ _1973_;
  assign _1978_ = b[27] & a[3];
  assign _1979_ = b[28] & a[2];
  assign _temp1263_ = _1979_ ^ _1978_;
  assign _1980_ = ~_temp1263_;
  assign _1981_ = b[29] & a[1];
  assign _1983_ = _1981_ ^ _1980_;
  assign _1984_ = ~_1983_;
  assign _1985_ = ~_1784_;
  assign _1986_ = _1783_ & _1782_;
  assign _temp1264_ = _1785_ & _1985_;
  assign _temp1265_ = _temp1264_ | _1986_;
  assign _1987_ = ~_temp1265_;
  assign _1988_ = _1987_ ^ _1984_;
  assign _1989_ = b[30] & a[0];
  assign _1990_ = _1989_ ^ _1988_;
  assign _1991_ = ~_1787_;
  assign _1992_ = _1788_ & _1991_;
  assign _1994_ = _1992_ ^ _1990_;
  assign _1995_ = _1994_ ^ _1977_;
  assign _1996_ = ~_1995_;
  assign _1997_ = _1996_ ^ _1946_;
  assign _1998_ = ~_1789_;
  assign _temp1266_ = _1780_ | _1777_;
  assign _1999_ = ~_temp1266_;
  assign _temp1267_ = _1998_ & _1781_;
  assign _temp1268_ = _temp1267_ | _1999_;
  assign _2000_ = ~_temp1268_;
  assign _2001_ = ~_2000_;
  assign _2002_ = _2001_ ^ _1997_;
  assign _2003_ = _2002_ ^ _1944_;
  assign _2005_ = _1746_ | _1743_;
  assign _temp1269_ = _1796_ | _1747_;
  assign _temp1270_ = _temp1269_ & _2005_;
  assign _2006_ = ~_temp1270_;
  assign _2007_ = _2006_ ^ _2003_;
  assign _2008_ = ~_1795_;
  assign _temp1271_ = _2008_ & _1791_;
  assign _2009_ = ~_temp1271_;
  assign _temp1272_ = _1790_ | _1751_;
  assign _temp1273_ = _temp1272_ & _2009_;
  assign _2010_ = ~_temp1273_;
  assign _2011_ = _2010_ ^ _2007_;
  assign _2012_ = ~_1798_;
  assign _2013_ = _1804_ | _1801_;
  assign _temp1274_ = _1800_ | _2012_;
  assign _temp1275_ = _temp1274_ & _2013_;
  assign _2014_ = ~_temp1275_;
  assign _2016_ = _2014_ ^ _2011_;
  assign _2017_ = _1809_ & _1805_;
  assign _2018_ = _2017_ ^ _2016_;
  assign _temp1276_ = _1811_ ^ _1810_;
  assign _2019_ = ~_temp1276_;
  assign _2020_ = _2019_ | _1608_;
  assign _2021_ = _1811_ & _1810_;
  assign _temp1277_ = _1813_ & _1812_;
  assign _temp1278_ = _temp1277_ | _2021_;
  assign _2022_ = ~_temp1278_;
  assign _temp1279_ = _2020_ | _1615_;
  assign _temp1280_ = _temp1279_ & _2022_;
  assign _2023_ = ~_temp1280_;
  assign q[30] = _2023_ ^ _2018_;
  assign _2024_ = a[31] & b[0];
  assign _2026_ = b[1] & a[30];
  assign _2027_ = _2026_ ^ _2024_;
  assign _2028_ = b[2] & a[29];
  assign _2029_ = _2028_ ^ _2027_;
  assign _2030_ = ~_1819_;
  assign _2031_ = _1817_ & _1816_;
  assign _temp1281_ = _1820_ & _2030_;
  assign _temp1282_ = _temp1281_ | _2031_;
  assign _2032_ = ~_temp1282_;
  assign _2033_ = _2032_ ^ _2029_;
  assign _temp1283_ = b[3] & a[28];
  assign _2034_ = ~_temp1283_;
  assign _2035_ = b[4] & a[27];
  assign _2036_ = _2035_ ^ _2034_;
  assign _2037_ = b[5] & a[26];
  assign _2038_ = _2037_ ^ _2036_;
  assign _2039_ = _2038_ ^ _2033_;
  assign _2040_ = _1824_ | _1821_;
  assign _2041_ = _1831_ | _1825_;
  assign _2042_ = _2041_ & _2040_;
  assign _2043_ = _2042_ ^ _2039_;
  assign _2044_ = ~_1828_;
  assign _2045_ = _1827_ & _1826_;
  assign _temp1284_ = _1830_ & _2044_;
  assign _temp1285_ = _temp1284_ | _2045_;
  assign _2048_ = ~_temp1285_;
  assign _temp1286_ = b[6] & a[25];
  assign _2049_ = ~_temp1286_;
  assign _2050_ = b[7] & a[24];
  assign _2051_ = _2050_ ^ _2049_;
  assign _2052_ = b[8] & a[23];
  assign _2053_ = _2052_ ^ _2051_;
  assign _2054_ = _2053_ ^ _2048_;
  assign _2055_ = ~_1843_;
  assign _2056_ = _1842_ & _1841_;
  assign _temp1287_ = _1844_ & _2055_;
  assign _temp1288_ = _temp1287_ | _2056_;
  assign _2057_ = ~_temp1288_;
  assign _2059_ = _2057_ ^ _2054_;
  assign _2060_ = _2059_ ^ _2043_;
  assign _temp1289_ = _1835_ | _1832_;
  assign _2061_ = ~_temp1289_;
  assign _temp1290_ = _1853_ & _1836_;
  assign _temp1291_ = _temp1290_ | _2061_;
  assign _2062_ = ~_temp1291_;
  assign _2063_ = _2062_ ^ _2060_;
  assign _2064_ = _1845_ | _1839_;
  assign _2065_ = _1850_ | _1846_;
  assign _2066_ = _2065_ & _2064_;
  assign _temp1292_ = b[9] & a[22];
  assign _2067_ = ~_temp1292_;
  assign _2068_ = b[10] & a[21];
  assign _2070_ = _2068_ ^ _2067_;
  assign _2071_ = b[11] & a[20];
  assign _2072_ = _2071_ ^ _2070_;
  assign _2073_ = ~_1864_;
  assign _2074_ = _1863_ & _1861_;
  assign _temp1293_ = _1865_ & _2073_;
  assign _temp1294_ = _temp1293_ | _2074_;
  assign _2075_ = ~_temp1294_;
  assign _2076_ = _2075_ ^ _2072_;
  assign _temp1295_ = b[12] & a[19];
  assign _2077_ = ~_temp1295_;
  assign _2078_ = b[13] & a[18];
  assign _2079_ = _2078_ ^ _2077_;
  assign _2081_ = b[14] & a[17];
  assign _2082_ = _2081_ ^ _2079_;
  assign _2083_ = _2082_ ^ _2076_;
  assign _2084_ = _2083_ ^ _2066_;
  assign _2085_ = _1869_ | _1866_;
  assign _2086_ = _1876_ | _1870_;
  assign _2087_ = _2086_ & _2085_;
  assign _2088_ = _2087_ ^ _2084_;
  assign _2089_ = _2088_ ^ _2063_;
  assign _2090_ = _1856_ & _1854_;
  assign _temp1296_ = _1886_ & _1857_;
  assign _temp1297_ = _temp1296_ | _2090_;
  assign _2092_ = ~_temp1297_;
  assign _2093_ = _2092_ ^ _2089_;
  assign _2094_ = _1878_ | _1860_;
  assign _2095_ = _1883_ | _1879_;
  assign _2096_ = _2095_ & _2094_;
  assign _2097_ = ~_1874_;
  assign _2098_ = _1872_ & _1871_;
  assign _temp1298_ = _1875_ & _2097_;
  assign _temp1299_ = _temp1298_ | _2098_;
  assign _2099_ = ~_temp1299_;
  assign _temp1300_ = b[15] & a[16];
  assign _2100_ = ~_temp1300_;
  assign _2101_ = b[16] & a[15];
  assign _2103_ = _2101_ ^ _2100_;
  assign _2104_ = b[17] & a[14];
  assign _2105_ = _2104_ ^ _2103_;
  assign _2106_ = _2105_ ^ _2099_;
  assign _2107_ = ~_1900_;
  assign _2108_ = _1899_ & _1898_;
  assign _temp1301_ = _1901_ & _2107_;
  assign _temp1302_ = _temp1301_ | _2108_;
  assign _2109_ = ~_temp1302_;
  assign _2110_ = _2109_ ^ _2106_;
  assign _2111_ = _1902_ | _1897_;
  assign _2112_ = _1907_ | _1903_;
  assign _2114_ = _2112_ & _2111_;
  assign _2115_ = _2114_ ^ _2110_;
  assign _temp1303_ = b[18] & a[13];
  assign _2116_ = ~_temp1303_;
  assign _2117_ = b[19] & a[12];
  assign _2118_ = _2117_ ^ _2116_;
  assign _2119_ = b[20] & a[11];
  assign _2120_ = _2119_ ^ _2118_;
  assign _2121_ = ~_1917_;
  assign _2122_ = _1915_ & _1914_;
  assign _temp1304_ = _1918_ & _2121_;
  assign _temp1305_ = _temp1304_ | _2122_;
  assign _2123_ = ~_temp1305_;
  assign _2125_ = _2123_ ^ _2120_;
  assign _temp1306_ = b[21] & a[10];
  assign _2126_ = ~_temp1306_;
  assign _2127_ = b[22] & a[9];
  assign _2128_ = _2127_ ^ _2126_;
  assign _2129_ = b[23] & a[8];
  assign _2130_ = _2129_ ^ _2128_;
  assign _2131_ = _2130_ ^ _2125_;
  assign _2132_ = _2131_ ^ _2115_;
  assign _2133_ = _2132_ ^ _2096_;
  assign _2134_ = _1912_ | _1909_;
  assign _2136_ = _1931_ | _1913_;
  assign _2137_ = _2136_ & _2134_;
  assign _2138_ = _2137_ ^ _2133_;
  assign _2139_ = _2138_ ^ _2093_;
  assign _2140_ = _1889_ & _1887_;
  assign _temp1307_ = _1940_ & _1890_;
  assign _temp1308_ = _temp1307_ | _2140_;
  assign _2141_ = ~_temp1308_;
  assign _2142_ = _2141_ ^ _2139_;
  assign _2143_ = _1933_ & _1893_;
  assign _temp1309_ = _1939_ & _1934_;
  assign _temp1310_ = _temp1309_ | _2143_;
  assign _2144_ = ~_temp1310_;
  assign _2145_ = _1922_ | _1919_;
  assign _2147_ = _1929_ | _1923_;
  assign _2148_ = _2147_ & _2145_;
  assign _2149_ = ~_1926_;
  assign _2150_ = _1925_ & _1924_;
  assign _temp1311_ = _1928_ & _2149_;
  assign _temp1312_ = _temp1311_ | _2150_;
  assign _2151_ = ~_temp1312_;
  assign _temp1313_ = a[7] & b[24];
  assign _2152_ = ~_temp1313_;
  assign _2153_ = b[25] & a[6];
  assign _2154_ = _2153_ ^ _2152_;
  assign _2155_ = b[26] & a[5];
  assign _2156_ = _2155_ ^ _2154_;
  assign _2158_ = _2156_ ^ _2151_;
  assign _2159_ = ~_1956_;
  assign _2160_ = _1955_ & _1954_;
  assign _temp1314_ = _1957_ & _2159_;
  assign _temp1315_ = _temp1314_ | _2160_;
  assign _2161_ = ~_temp1315_;
  assign _2162_ = _2161_ ^ _2158_;
  assign _2163_ = _2162_ ^ _2148_;
  assign _2164_ = _1958_ | _1953_;
  assign _2165_ = _1964_ | _1959_;
  assign _2166_ = _2165_ & _2164_;
  assign _2167_ = _2166_ ^ _2163_;
  assign _2169_ = _1966_ | _1950_;
  assign _2170_ = _1972_ | _1967_;
  assign _2171_ = _2170_ & _2169_;
  assign _2172_ = _2171_ ^ _2167_;
  assign _temp1316_ = b[27] & a[4];
  assign _2173_ = ~_temp1316_;
  assign _2174_ = b[28] & a[3];
  assign _2175_ = _2174_ ^ _2173_;
  assign _2176_ = b[29] & a[2];
  assign _2177_ = _2176_ ^ _2175_;
  assign _2178_ = ~_1980_;
  assign _2180_ = _1979_ & _1978_;
  assign _temp1317_ = _1981_ & _2178_;
  assign _temp1318_ = _temp1317_ | _2180_;
  assign _2181_ = ~_temp1318_;
  assign _2182_ = _2181_ ^ _2177_;
  assign _2183_ = b[30] & a[1];
  assign _2184_ = _2183_ ^ _2182_;
  assign _2185_ = ~_1988_;
  assign _temp1319_ = _1987_ | _1983_;
  assign _2186_ = ~_temp1319_;
  assign _temp1320_ = _1989_ & _2185_;
  assign _temp1321_ = _temp1320_ | _2186_;
  assign _2187_ = ~_temp1321_;
  assign _2188_ = _2187_ ^ _2184_;
  assign _2189_ = b[31] & a[0];
  assign _2191_ = _2189_ ^ _2188_;
  assign _2192_ = _2191_ ^ _2172_;
  assign _2193_ = _2192_ ^ _2144_;
  assign _2194_ = ~_1994_;
  assign _temp1322_ = _1976_ | _1973_;
  assign _2195_ = ~_temp1322_;
  assign _temp1323_ = _2194_ & _1977_;
  assign _temp1324_ = _temp1323_ | _2195_;
  assign _2196_ = ~_temp1324_;
  assign _2197_ = _2196_ ^ _2193_;
  assign _2198_ = _2197_ ^ _2142_;
  assign _2199_ = _1943_ & _1941_;
  assign _temp1325_ = _2002_ & _1944_;
  assign _temp1326_ = _temp1325_ | _2199_;
  assign _2200_ = ~_temp1326_;
  assign _2202_ = _2200_ ^ _2198_;
  assign _2203_ = _1996_ & _1946_;
  assign _temp1327_ = _2001_ & _1997_;
  assign _temp1328_ = _temp1327_ | _2203_;
  assign _2204_ = ~_temp1328_;
  assign _2205_ = _2204_ ^ _2202_;
  assign _2206_ = _2006_ & _2003_;
  assign _temp1329_ = _2010_ & _2007_;
  assign _temp1330_ = _temp1329_ | _2206_;
  assign _2207_ = ~_temp1330_;
  assign _2208_ = _2207_ ^ _2205_;
  assign _2209_ = ~_1990_;
  assign _2210_ = _1992_ & _2209_;
  assign _2211_ = _2210_ ^ _2208_;
  assign _2213_ = _2014_ & _2011_;
  assign _2214_ = _2213_ ^ _2211_;
  assign _2215_ = _2017_ & _2016_;
  assign _temp1331_ = _2023_ & _2018_;
  assign _temp1332_ = _temp1331_ | _2215_;
  assign _2216_ = ~_temp1332_;
  assign q[31] = _2216_ ^ _2214_;
endmodule
