module or_gate(q, a, b);
    output q;
    input a, b;
    assign q = a | b;
endmodule
